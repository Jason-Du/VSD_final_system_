# 
#              Synchronous Dual Port SRAM Compiler 
# 
#                    UMC 0.18um Generic Logic Process 
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2009 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http://www.faraday-tech.com/
#   
#       Module Name      : layer1_sram
#       Words            : 912
#       Bits             : 128
#       Byte-Write       : 1
#       Aspect Ratio     : 1
#       Output Loading   : 0.5  (pf)
#       Data Slew        : 2.0  (ns)
#       CK Slew          : 2.0  (ns)
#       Power Ring Width : 2  (um)
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSA0M_A
#       Memaker          : 200901.2.1
#       Date             : 2021/01/15 13:25:24
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO layer1_sram
CLASS BLOCK ;
FOREIGN layer1_sram 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 3596.000 BY 501.760 ;
SYMMETRY x y r90 ;
SITE core ;
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal5 ;
  RECT 3594.880 489.780 3596.000 493.020 ;
  LAYER metal4 ;
  RECT 3594.880 489.780 3596.000 493.020 ;
  LAYER metal3 ;
  RECT 3594.880 489.780 3596.000 493.020 ;
  LAYER metal2 ;
  RECT 3594.880 489.780 3596.000 493.020 ;
  LAYER metal1 ;
  RECT 3594.880 489.780 3596.000 493.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 481.940 3596.000 485.180 ;
  LAYER metal4 ;
  RECT 3594.880 481.940 3596.000 485.180 ;
  LAYER metal3 ;
  RECT 3594.880 481.940 3596.000 485.180 ;
  LAYER metal2 ;
  RECT 3594.880 481.940 3596.000 485.180 ;
  LAYER metal1 ;
  RECT 3594.880 481.940 3596.000 485.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 442.740 3596.000 445.980 ;
  LAYER metal4 ;
  RECT 3594.880 442.740 3596.000 445.980 ;
  LAYER metal3 ;
  RECT 3594.880 442.740 3596.000 445.980 ;
  LAYER metal2 ;
  RECT 3594.880 442.740 3596.000 445.980 ;
  LAYER metal1 ;
  RECT 3594.880 442.740 3596.000 445.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 434.900 3596.000 438.140 ;
  LAYER metal4 ;
  RECT 3594.880 434.900 3596.000 438.140 ;
  LAYER metal3 ;
  RECT 3594.880 434.900 3596.000 438.140 ;
  LAYER metal2 ;
  RECT 3594.880 434.900 3596.000 438.140 ;
  LAYER metal1 ;
  RECT 3594.880 434.900 3596.000 438.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 427.060 3596.000 430.300 ;
  LAYER metal4 ;
  RECT 3594.880 427.060 3596.000 430.300 ;
  LAYER metal3 ;
  RECT 3594.880 427.060 3596.000 430.300 ;
  LAYER metal2 ;
  RECT 3594.880 427.060 3596.000 430.300 ;
  LAYER metal1 ;
  RECT 3594.880 427.060 3596.000 430.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 419.220 3596.000 422.460 ;
  LAYER metal4 ;
  RECT 3594.880 419.220 3596.000 422.460 ;
  LAYER metal3 ;
  RECT 3594.880 419.220 3596.000 422.460 ;
  LAYER metal2 ;
  RECT 3594.880 419.220 3596.000 422.460 ;
  LAYER metal1 ;
  RECT 3594.880 419.220 3596.000 422.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 411.380 3596.000 414.620 ;
  LAYER metal4 ;
  RECT 3594.880 411.380 3596.000 414.620 ;
  LAYER metal3 ;
  RECT 3594.880 411.380 3596.000 414.620 ;
  LAYER metal2 ;
  RECT 3594.880 411.380 3596.000 414.620 ;
  LAYER metal1 ;
  RECT 3594.880 411.380 3596.000 414.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 403.540 3596.000 406.780 ;
  LAYER metal4 ;
  RECT 3594.880 403.540 3596.000 406.780 ;
  LAYER metal3 ;
  RECT 3594.880 403.540 3596.000 406.780 ;
  LAYER metal2 ;
  RECT 3594.880 403.540 3596.000 406.780 ;
  LAYER metal1 ;
  RECT 3594.880 403.540 3596.000 406.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 364.340 3596.000 367.580 ;
  LAYER metal4 ;
  RECT 3594.880 364.340 3596.000 367.580 ;
  LAYER metal3 ;
  RECT 3594.880 364.340 3596.000 367.580 ;
  LAYER metal2 ;
  RECT 3594.880 364.340 3596.000 367.580 ;
  LAYER metal1 ;
  RECT 3594.880 364.340 3596.000 367.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 356.500 3596.000 359.740 ;
  LAYER metal4 ;
  RECT 3594.880 356.500 3596.000 359.740 ;
  LAYER metal3 ;
  RECT 3594.880 356.500 3596.000 359.740 ;
  LAYER metal2 ;
  RECT 3594.880 356.500 3596.000 359.740 ;
  LAYER metal1 ;
  RECT 3594.880 356.500 3596.000 359.740 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 348.660 3596.000 351.900 ;
  LAYER metal4 ;
  RECT 3594.880 348.660 3596.000 351.900 ;
  LAYER metal3 ;
  RECT 3594.880 348.660 3596.000 351.900 ;
  LAYER metal2 ;
  RECT 3594.880 348.660 3596.000 351.900 ;
  LAYER metal1 ;
  RECT 3594.880 348.660 3596.000 351.900 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 340.820 3596.000 344.060 ;
  LAYER metal4 ;
  RECT 3594.880 340.820 3596.000 344.060 ;
  LAYER metal3 ;
  RECT 3594.880 340.820 3596.000 344.060 ;
  LAYER metal2 ;
  RECT 3594.880 340.820 3596.000 344.060 ;
  LAYER metal1 ;
  RECT 3594.880 340.820 3596.000 344.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 332.980 3596.000 336.220 ;
  LAYER metal4 ;
  RECT 3594.880 332.980 3596.000 336.220 ;
  LAYER metal3 ;
  RECT 3594.880 332.980 3596.000 336.220 ;
  LAYER metal2 ;
  RECT 3594.880 332.980 3596.000 336.220 ;
  LAYER metal1 ;
  RECT 3594.880 332.980 3596.000 336.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 325.140 3596.000 328.380 ;
  LAYER metal4 ;
  RECT 3594.880 325.140 3596.000 328.380 ;
  LAYER metal3 ;
  RECT 3594.880 325.140 3596.000 328.380 ;
  LAYER metal2 ;
  RECT 3594.880 325.140 3596.000 328.380 ;
  LAYER metal1 ;
  RECT 3594.880 325.140 3596.000 328.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 285.940 3596.000 289.180 ;
  LAYER metal4 ;
  RECT 3594.880 285.940 3596.000 289.180 ;
  LAYER metal3 ;
  RECT 3594.880 285.940 3596.000 289.180 ;
  LAYER metal2 ;
  RECT 3594.880 285.940 3596.000 289.180 ;
  LAYER metal1 ;
  RECT 3594.880 285.940 3596.000 289.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 278.100 3596.000 281.340 ;
  LAYER metal4 ;
  RECT 3594.880 278.100 3596.000 281.340 ;
  LAYER metal3 ;
  RECT 3594.880 278.100 3596.000 281.340 ;
  LAYER metal2 ;
  RECT 3594.880 278.100 3596.000 281.340 ;
  LAYER metal1 ;
  RECT 3594.880 278.100 3596.000 281.340 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 270.260 3596.000 273.500 ;
  LAYER metal4 ;
  RECT 3594.880 270.260 3596.000 273.500 ;
  LAYER metal3 ;
  RECT 3594.880 270.260 3596.000 273.500 ;
  LAYER metal2 ;
  RECT 3594.880 270.260 3596.000 273.500 ;
  LAYER metal1 ;
  RECT 3594.880 270.260 3596.000 273.500 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 262.420 3596.000 265.660 ;
  LAYER metal4 ;
  RECT 3594.880 262.420 3596.000 265.660 ;
  LAYER metal3 ;
  RECT 3594.880 262.420 3596.000 265.660 ;
  LAYER metal2 ;
  RECT 3594.880 262.420 3596.000 265.660 ;
  LAYER metal1 ;
  RECT 3594.880 262.420 3596.000 265.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 254.580 3596.000 257.820 ;
  LAYER metal4 ;
  RECT 3594.880 254.580 3596.000 257.820 ;
  LAYER metal3 ;
  RECT 3594.880 254.580 3596.000 257.820 ;
  LAYER metal2 ;
  RECT 3594.880 254.580 3596.000 257.820 ;
  LAYER metal1 ;
  RECT 3594.880 254.580 3596.000 257.820 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 246.740 3596.000 249.980 ;
  LAYER metal4 ;
  RECT 3594.880 246.740 3596.000 249.980 ;
  LAYER metal3 ;
  RECT 3594.880 246.740 3596.000 249.980 ;
  LAYER metal2 ;
  RECT 3594.880 246.740 3596.000 249.980 ;
  LAYER metal1 ;
  RECT 3594.880 246.740 3596.000 249.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 207.540 3596.000 210.780 ;
  LAYER metal4 ;
  RECT 3594.880 207.540 3596.000 210.780 ;
  LAYER metal3 ;
  RECT 3594.880 207.540 3596.000 210.780 ;
  LAYER metal2 ;
  RECT 3594.880 207.540 3596.000 210.780 ;
  LAYER metal1 ;
  RECT 3594.880 207.540 3596.000 210.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 199.700 3596.000 202.940 ;
  LAYER metal4 ;
  RECT 3594.880 199.700 3596.000 202.940 ;
  LAYER metal3 ;
  RECT 3594.880 199.700 3596.000 202.940 ;
  LAYER metal2 ;
  RECT 3594.880 199.700 3596.000 202.940 ;
  LAYER metal1 ;
  RECT 3594.880 199.700 3596.000 202.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 191.860 3596.000 195.100 ;
  LAYER metal4 ;
  RECT 3594.880 191.860 3596.000 195.100 ;
  LAYER metal3 ;
  RECT 3594.880 191.860 3596.000 195.100 ;
  LAYER metal2 ;
  RECT 3594.880 191.860 3596.000 195.100 ;
  LAYER metal1 ;
  RECT 3594.880 191.860 3596.000 195.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 184.020 3596.000 187.260 ;
  LAYER metal4 ;
  RECT 3594.880 184.020 3596.000 187.260 ;
  LAYER metal3 ;
  RECT 3594.880 184.020 3596.000 187.260 ;
  LAYER metal2 ;
  RECT 3594.880 184.020 3596.000 187.260 ;
  LAYER metal1 ;
  RECT 3594.880 184.020 3596.000 187.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 176.180 3596.000 179.420 ;
  LAYER metal4 ;
  RECT 3594.880 176.180 3596.000 179.420 ;
  LAYER metal3 ;
  RECT 3594.880 176.180 3596.000 179.420 ;
  LAYER metal2 ;
  RECT 3594.880 176.180 3596.000 179.420 ;
  LAYER metal1 ;
  RECT 3594.880 176.180 3596.000 179.420 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 168.340 3596.000 171.580 ;
  LAYER metal4 ;
  RECT 3594.880 168.340 3596.000 171.580 ;
  LAYER metal3 ;
  RECT 3594.880 168.340 3596.000 171.580 ;
  LAYER metal2 ;
  RECT 3594.880 168.340 3596.000 171.580 ;
  LAYER metal1 ;
  RECT 3594.880 168.340 3596.000 171.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 129.140 3596.000 132.380 ;
  LAYER metal4 ;
  RECT 3594.880 129.140 3596.000 132.380 ;
  LAYER metal3 ;
  RECT 3594.880 129.140 3596.000 132.380 ;
  LAYER metal2 ;
  RECT 3594.880 129.140 3596.000 132.380 ;
  LAYER metal1 ;
  RECT 3594.880 129.140 3596.000 132.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 121.300 3596.000 124.540 ;
  LAYER metal4 ;
  RECT 3594.880 121.300 3596.000 124.540 ;
  LAYER metal3 ;
  RECT 3594.880 121.300 3596.000 124.540 ;
  LAYER metal2 ;
  RECT 3594.880 121.300 3596.000 124.540 ;
  LAYER metal1 ;
  RECT 3594.880 121.300 3596.000 124.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 113.460 3596.000 116.700 ;
  LAYER metal4 ;
  RECT 3594.880 113.460 3596.000 116.700 ;
  LAYER metal3 ;
  RECT 3594.880 113.460 3596.000 116.700 ;
  LAYER metal2 ;
  RECT 3594.880 113.460 3596.000 116.700 ;
  LAYER metal1 ;
  RECT 3594.880 113.460 3596.000 116.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 105.620 3596.000 108.860 ;
  LAYER metal4 ;
  RECT 3594.880 105.620 3596.000 108.860 ;
  LAYER metal3 ;
  RECT 3594.880 105.620 3596.000 108.860 ;
  LAYER metal2 ;
  RECT 3594.880 105.620 3596.000 108.860 ;
  LAYER metal1 ;
  RECT 3594.880 105.620 3596.000 108.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 97.780 3596.000 101.020 ;
  LAYER metal4 ;
  RECT 3594.880 97.780 3596.000 101.020 ;
  LAYER metal3 ;
  RECT 3594.880 97.780 3596.000 101.020 ;
  LAYER metal2 ;
  RECT 3594.880 97.780 3596.000 101.020 ;
  LAYER metal1 ;
  RECT 3594.880 97.780 3596.000 101.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 89.940 3596.000 93.180 ;
  LAYER metal4 ;
  RECT 3594.880 89.940 3596.000 93.180 ;
  LAYER metal3 ;
  RECT 3594.880 89.940 3596.000 93.180 ;
  LAYER metal2 ;
  RECT 3594.880 89.940 3596.000 93.180 ;
  LAYER metal1 ;
  RECT 3594.880 89.940 3596.000 93.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 50.740 3596.000 53.980 ;
  LAYER metal4 ;
  RECT 3594.880 50.740 3596.000 53.980 ;
  LAYER metal3 ;
  RECT 3594.880 50.740 3596.000 53.980 ;
  LAYER metal2 ;
  RECT 3594.880 50.740 3596.000 53.980 ;
  LAYER metal1 ;
  RECT 3594.880 50.740 3596.000 53.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 42.900 3596.000 46.140 ;
  LAYER metal4 ;
  RECT 3594.880 42.900 3596.000 46.140 ;
  LAYER metal3 ;
  RECT 3594.880 42.900 3596.000 46.140 ;
  LAYER metal2 ;
  RECT 3594.880 42.900 3596.000 46.140 ;
  LAYER metal1 ;
  RECT 3594.880 42.900 3596.000 46.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 35.060 3596.000 38.300 ;
  LAYER metal4 ;
  RECT 3594.880 35.060 3596.000 38.300 ;
  LAYER metal3 ;
  RECT 3594.880 35.060 3596.000 38.300 ;
  LAYER metal2 ;
  RECT 3594.880 35.060 3596.000 38.300 ;
  LAYER metal1 ;
  RECT 3594.880 35.060 3596.000 38.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 27.220 3596.000 30.460 ;
  LAYER metal4 ;
  RECT 3594.880 27.220 3596.000 30.460 ;
  LAYER metal3 ;
  RECT 3594.880 27.220 3596.000 30.460 ;
  LAYER metal2 ;
  RECT 3594.880 27.220 3596.000 30.460 ;
  LAYER metal1 ;
  RECT 3594.880 27.220 3596.000 30.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 19.380 3596.000 22.620 ;
  LAYER metal4 ;
  RECT 3594.880 19.380 3596.000 22.620 ;
  LAYER metal3 ;
  RECT 3594.880 19.380 3596.000 22.620 ;
  LAYER metal2 ;
  RECT 3594.880 19.380 3596.000 22.620 ;
  LAYER metal1 ;
  RECT 3594.880 19.380 3596.000 22.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 11.540 3596.000 14.780 ;
  LAYER metal4 ;
  RECT 3594.880 11.540 3596.000 14.780 ;
  LAYER metal3 ;
  RECT 3594.880 11.540 3596.000 14.780 ;
  LAYER metal2 ;
  RECT 3594.880 11.540 3596.000 14.780 ;
  LAYER metal1 ;
  RECT 3594.880 11.540 3596.000 14.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 489.780 1.120 493.020 ;
  LAYER metal4 ;
  RECT 0.000 489.780 1.120 493.020 ;
  LAYER metal3 ;
  RECT 0.000 489.780 1.120 493.020 ;
  LAYER metal2 ;
  RECT 0.000 489.780 1.120 493.020 ;
  LAYER metal1 ;
  RECT 0.000 489.780 1.120 493.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 481.940 1.120 485.180 ;
  LAYER metal4 ;
  RECT 0.000 481.940 1.120 485.180 ;
  LAYER metal3 ;
  RECT 0.000 481.940 1.120 485.180 ;
  LAYER metal2 ;
  RECT 0.000 481.940 1.120 485.180 ;
  LAYER metal1 ;
  RECT 0.000 481.940 1.120 485.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 442.740 1.120 445.980 ;
  LAYER metal4 ;
  RECT 0.000 442.740 1.120 445.980 ;
  LAYER metal3 ;
  RECT 0.000 442.740 1.120 445.980 ;
  LAYER metal2 ;
  RECT 0.000 442.740 1.120 445.980 ;
  LAYER metal1 ;
  RECT 0.000 442.740 1.120 445.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 434.900 1.120 438.140 ;
  LAYER metal4 ;
  RECT 0.000 434.900 1.120 438.140 ;
  LAYER metal3 ;
  RECT 0.000 434.900 1.120 438.140 ;
  LAYER metal2 ;
  RECT 0.000 434.900 1.120 438.140 ;
  LAYER metal1 ;
  RECT 0.000 434.900 1.120 438.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 427.060 1.120 430.300 ;
  LAYER metal4 ;
  RECT 0.000 427.060 1.120 430.300 ;
  LAYER metal3 ;
  RECT 0.000 427.060 1.120 430.300 ;
  LAYER metal2 ;
  RECT 0.000 427.060 1.120 430.300 ;
  LAYER metal1 ;
  RECT 0.000 427.060 1.120 430.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 419.220 1.120 422.460 ;
  LAYER metal4 ;
  RECT 0.000 419.220 1.120 422.460 ;
  LAYER metal3 ;
  RECT 0.000 419.220 1.120 422.460 ;
  LAYER metal2 ;
  RECT 0.000 419.220 1.120 422.460 ;
  LAYER metal1 ;
  RECT 0.000 419.220 1.120 422.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 411.380 1.120 414.620 ;
  LAYER metal4 ;
  RECT 0.000 411.380 1.120 414.620 ;
  LAYER metal3 ;
  RECT 0.000 411.380 1.120 414.620 ;
  LAYER metal2 ;
  RECT 0.000 411.380 1.120 414.620 ;
  LAYER metal1 ;
  RECT 0.000 411.380 1.120 414.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 403.540 1.120 406.780 ;
  LAYER metal4 ;
  RECT 0.000 403.540 1.120 406.780 ;
  LAYER metal3 ;
  RECT 0.000 403.540 1.120 406.780 ;
  LAYER metal2 ;
  RECT 0.000 403.540 1.120 406.780 ;
  LAYER metal1 ;
  RECT 0.000 403.540 1.120 406.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 364.340 1.120 367.580 ;
  LAYER metal4 ;
  RECT 0.000 364.340 1.120 367.580 ;
  LAYER metal3 ;
  RECT 0.000 364.340 1.120 367.580 ;
  LAYER metal2 ;
  RECT 0.000 364.340 1.120 367.580 ;
  LAYER metal1 ;
  RECT 0.000 364.340 1.120 367.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 356.500 1.120 359.740 ;
  LAYER metal4 ;
  RECT 0.000 356.500 1.120 359.740 ;
  LAYER metal3 ;
  RECT 0.000 356.500 1.120 359.740 ;
  LAYER metal2 ;
  RECT 0.000 356.500 1.120 359.740 ;
  LAYER metal1 ;
  RECT 0.000 356.500 1.120 359.740 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 348.660 1.120 351.900 ;
  LAYER metal4 ;
  RECT 0.000 348.660 1.120 351.900 ;
  LAYER metal3 ;
  RECT 0.000 348.660 1.120 351.900 ;
  LAYER metal2 ;
  RECT 0.000 348.660 1.120 351.900 ;
  LAYER metal1 ;
  RECT 0.000 348.660 1.120 351.900 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 340.820 1.120 344.060 ;
  LAYER metal4 ;
  RECT 0.000 340.820 1.120 344.060 ;
  LAYER metal3 ;
  RECT 0.000 340.820 1.120 344.060 ;
  LAYER metal2 ;
  RECT 0.000 340.820 1.120 344.060 ;
  LAYER metal1 ;
  RECT 0.000 340.820 1.120 344.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 332.980 1.120 336.220 ;
  LAYER metal4 ;
  RECT 0.000 332.980 1.120 336.220 ;
  LAYER metal3 ;
  RECT 0.000 332.980 1.120 336.220 ;
  LAYER metal2 ;
  RECT 0.000 332.980 1.120 336.220 ;
  LAYER metal1 ;
  RECT 0.000 332.980 1.120 336.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 325.140 1.120 328.380 ;
  LAYER metal4 ;
  RECT 0.000 325.140 1.120 328.380 ;
  LAYER metal3 ;
  RECT 0.000 325.140 1.120 328.380 ;
  LAYER metal2 ;
  RECT 0.000 325.140 1.120 328.380 ;
  LAYER metal1 ;
  RECT 0.000 325.140 1.120 328.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 285.940 1.120 289.180 ;
  LAYER metal4 ;
  RECT 0.000 285.940 1.120 289.180 ;
  LAYER metal3 ;
  RECT 0.000 285.940 1.120 289.180 ;
  LAYER metal2 ;
  RECT 0.000 285.940 1.120 289.180 ;
  LAYER metal1 ;
  RECT 0.000 285.940 1.120 289.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 278.100 1.120 281.340 ;
  LAYER metal4 ;
  RECT 0.000 278.100 1.120 281.340 ;
  LAYER metal3 ;
  RECT 0.000 278.100 1.120 281.340 ;
  LAYER metal2 ;
  RECT 0.000 278.100 1.120 281.340 ;
  LAYER metal1 ;
  RECT 0.000 278.100 1.120 281.340 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 270.260 1.120 273.500 ;
  LAYER metal4 ;
  RECT 0.000 270.260 1.120 273.500 ;
  LAYER metal3 ;
  RECT 0.000 270.260 1.120 273.500 ;
  LAYER metal2 ;
  RECT 0.000 270.260 1.120 273.500 ;
  LAYER metal1 ;
  RECT 0.000 270.260 1.120 273.500 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 262.420 1.120 265.660 ;
  LAYER metal4 ;
  RECT 0.000 262.420 1.120 265.660 ;
  LAYER metal3 ;
  RECT 0.000 262.420 1.120 265.660 ;
  LAYER metal2 ;
  RECT 0.000 262.420 1.120 265.660 ;
  LAYER metal1 ;
  RECT 0.000 262.420 1.120 265.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 254.580 1.120 257.820 ;
  LAYER metal4 ;
  RECT 0.000 254.580 1.120 257.820 ;
  LAYER metal3 ;
  RECT 0.000 254.580 1.120 257.820 ;
  LAYER metal2 ;
  RECT 0.000 254.580 1.120 257.820 ;
  LAYER metal1 ;
  RECT 0.000 254.580 1.120 257.820 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 246.740 1.120 249.980 ;
  LAYER metal4 ;
  RECT 0.000 246.740 1.120 249.980 ;
  LAYER metal3 ;
  RECT 0.000 246.740 1.120 249.980 ;
  LAYER metal2 ;
  RECT 0.000 246.740 1.120 249.980 ;
  LAYER metal1 ;
  RECT 0.000 246.740 1.120 249.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 207.540 1.120 210.780 ;
  LAYER metal4 ;
  RECT 0.000 207.540 1.120 210.780 ;
  LAYER metal3 ;
  RECT 0.000 207.540 1.120 210.780 ;
  LAYER metal2 ;
  RECT 0.000 207.540 1.120 210.780 ;
  LAYER metal1 ;
  RECT 0.000 207.540 1.120 210.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 199.700 1.120 202.940 ;
  LAYER metal4 ;
  RECT 0.000 199.700 1.120 202.940 ;
  LAYER metal3 ;
  RECT 0.000 199.700 1.120 202.940 ;
  LAYER metal2 ;
  RECT 0.000 199.700 1.120 202.940 ;
  LAYER metal1 ;
  RECT 0.000 199.700 1.120 202.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 191.860 1.120 195.100 ;
  LAYER metal4 ;
  RECT 0.000 191.860 1.120 195.100 ;
  LAYER metal3 ;
  RECT 0.000 191.860 1.120 195.100 ;
  LAYER metal2 ;
  RECT 0.000 191.860 1.120 195.100 ;
  LAYER metal1 ;
  RECT 0.000 191.860 1.120 195.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 184.020 1.120 187.260 ;
  LAYER metal4 ;
  RECT 0.000 184.020 1.120 187.260 ;
  LAYER metal3 ;
  RECT 0.000 184.020 1.120 187.260 ;
  LAYER metal2 ;
  RECT 0.000 184.020 1.120 187.260 ;
  LAYER metal1 ;
  RECT 0.000 184.020 1.120 187.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 176.180 1.120 179.420 ;
  LAYER metal4 ;
  RECT 0.000 176.180 1.120 179.420 ;
  LAYER metal3 ;
  RECT 0.000 176.180 1.120 179.420 ;
  LAYER metal2 ;
  RECT 0.000 176.180 1.120 179.420 ;
  LAYER metal1 ;
  RECT 0.000 176.180 1.120 179.420 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 168.340 1.120 171.580 ;
  LAYER metal4 ;
  RECT 0.000 168.340 1.120 171.580 ;
  LAYER metal3 ;
  RECT 0.000 168.340 1.120 171.580 ;
  LAYER metal2 ;
  RECT 0.000 168.340 1.120 171.580 ;
  LAYER metal1 ;
  RECT 0.000 168.340 1.120 171.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 129.140 1.120 132.380 ;
  LAYER metal4 ;
  RECT 0.000 129.140 1.120 132.380 ;
  LAYER metal3 ;
  RECT 0.000 129.140 1.120 132.380 ;
  LAYER metal2 ;
  RECT 0.000 129.140 1.120 132.380 ;
  LAYER metal1 ;
  RECT 0.000 129.140 1.120 132.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 121.300 1.120 124.540 ;
  LAYER metal4 ;
  RECT 0.000 121.300 1.120 124.540 ;
  LAYER metal3 ;
  RECT 0.000 121.300 1.120 124.540 ;
  LAYER metal2 ;
  RECT 0.000 121.300 1.120 124.540 ;
  LAYER metal1 ;
  RECT 0.000 121.300 1.120 124.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 113.460 1.120 116.700 ;
  LAYER metal4 ;
  RECT 0.000 113.460 1.120 116.700 ;
  LAYER metal3 ;
  RECT 0.000 113.460 1.120 116.700 ;
  LAYER metal2 ;
  RECT 0.000 113.460 1.120 116.700 ;
  LAYER metal1 ;
  RECT 0.000 113.460 1.120 116.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 105.620 1.120 108.860 ;
  LAYER metal4 ;
  RECT 0.000 105.620 1.120 108.860 ;
  LAYER metal3 ;
  RECT 0.000 105.620 1.120 108.860 ;
  LAYER metal2 ;
  RECT 0.000 105.620 1.120 108.860 ;
  LAYER metal1 ;
  RECT 0.000 105.620 1.120 108.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 97.780 1.120 101.020 ;
  LAYER metal4 ;
  RECT 0.000 97.780 1.120 101.020 ;
  LAYER metal3 ;
  RECT 0.000 97.780 1.120 101.020 ;
  LAYER metal2 ;
  RECT 0.000 97.780 1.120 101.020 ;
  LAYER metal1 ;
  RECT 0.000 97.780 1.120 101.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 89.940 1.120 93.180 ;
  LAYER metal4 ;
  RECT 0.000 89.940 1.120 93.180 ;
  LAYER metal3 ;
  RECT 0.000 89.940 1.120 93.180 ;
  LAYER metal2 ;
  RECT 0.000 89.940 1.120 93.180 ;
  LAYER metal1 ;
  RECT 0.000 89.940 1.120 93.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 50.740 1.120 53.980 ;
  LAYER metal4 ;
  RECT 0.000 50.740 1.120 53.980 ;
  LAYER metal3 ;
  RECT 0.000 50.740 1.120 53.980 ;
  LAYER metal2 ;
  RECT 0.000 50.740 1.120 53.980 ;
  LAYER metal1 ;
  RECT 0.000 50.740 1.120 53.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 42.900 1.120 46.140 ;
  LAYER metal4 ;
  RECT 0.000 42.900 1.120 46.140 ;
  LAYER metal3 ;
  RECT 0.000 42.900 1.120 46.140 ;
  LAYER metal2 ;
  RECT 0.000 42.900 1.120 46.140 ;
  LAYER metal1 ;
  RECT 0.000 42.900 1.120 46.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 35.060 1.120 38.300 ;
  LAYER metal4 ;
  RECT 0.000 35.060 1.120 38.300 ;
  LAYER metal3 ;
  RECT 0.000 35.060 1.120 38.300 ;
  LAYER metal2 ;
  RECT 0.000 35.060 1.120 38.300 ;
  LAYER metal1 ;
  RECT 0.000 35.060 1.120 38.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 27.220 1.120 30.460 ;
  LAYER metal4 ;
  RECT 0.000 27.220 1.120 30.460 ;
  LAYER metal3 ;
  RECT 0.000 27.220 1.120 30.460 ;
  LAYER metal2 ;
  RECT 0.000 27.220 1.120 30.460 ;
  LAYER metal1 ;
  RECT 0.000 27.220 1.120 30.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 19.380 1.120 22.620 ;
  LAYER metal4 ;
  RECT 0.000 19.380 1.120 22.620 ;
  LAYER metal3 ;
  RECT 0.000 19.380 1.120 22.620 ;
  LAYER metal2 ;
  RECT 0.000 19.380 1.120 22.620 ;
  LAYER metal1 ;
  RECT 0.000 19.380 1.120 22.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 11.540 1.120 14.780 ;
  LAYER metal4 ;
  RECT 0.000 11.540 1.120 14.780 ;
  LAYER metal3 ;
  RECT 0.000 11.540 1.120 14.780 ;
  LAYER metal2 ;
  RECT 0.000 11.540 1.120 14.780 ;
  LAYER metal1 ;
  RECT 0.000 11.540 1.120 14.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3579.660 500.640 3583.200 501.760 ;
  LAYER metal4 ;
  RECT 3579.660 500.640 3583.200 501.760 ;
  LAYER metal3 ;
  RECT 3579.660 500.640 3583.200 501.760 ;
  LAYER metal2 ;
  RECT 3579.660 500.640 3583.200 501.760 ;
  LAYER metal1 ;
  RECT 3579.660 500.640 3583.200 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3566.020 500.640 3569.560 501.760 ;
  LAYER metal4 ;
  RECT 3566.020 500.640 3569.560 501.760 ;
  LAYER metal3 ;
  RECT 3566.020 500.640 3569.560 501.760 ;
  LAYER metal2 ;
  RECT 3566.020 500.640 3569.560 501.760 ;
  LAYER metal1 ;
  RECT 3566.020 500.640 3569.560 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3553.000 500.640 3556.540 501.760 ;
  LAYER metal4 ;
  RECT 3553.000 500.640 3556.540 501.760 ;
  LAYER metal3 ;
  RECT 3553.000 500.640 3556.540 501.760 ;
  LAYER metal2 ;
  RECT 3553.000 500.640 3556.540 501.760 ;
  LAYER metal1 ;
  RECT 3553.000 500.640 3556.540 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3539.360 500.640 3542.900 501.760 ;
  LAYER metal4 ;
  RECT 3539.360 500.640 3542.900 501.760 ;
  LAYER metal3 ;
  RECT 3539.360 500.640 3542.900 501.760 ;
  LAYER metal2 ;
  RECT 3539.360 500.640 3542.900 501.760 ;
  LAYER metal1 ;
  RECT 3539.360 500.640 3542.900 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3525.720 500.640 3529.260 501.760 ;
  LAYER metal4 ;
  RECT 3525.720 500.640 3529.260 501.760 ;
  LAYER metal3 ;
  RECT 3525.720 500.640 3529.260 501.760 ;
  LAYER metal2 ;
  RECT 3525.720 500.640 3529.260 501.760 ;
  LAYER metal1 ;
  RECT 3525.720 500.640 3529.260 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3458.760 500.640 3462.300 501.760 ;
  LAYER metal4 ;
  RECT 3458.760 500.640 3462.300 501.760 ;
  LAYER metal3 ;
  RECT 3458.760 500.640 3462.300 501.760 ;
  LAYER metal2 ;
  RECT 3458.760 500.640 3462.300 501.760 ;
  LAYER metal1 ;
  RECT 3458.760 500.640 3462.300 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3445.120 500.640 3448.660 501.760 ;
  LAYER metal4 ;
  RECT 3445.120 500.640 3448.660 501.760 ;
  LAYER metal3 ;
  RECT 3445.120 500.640 3448.660 501.760 ;
  LAYER metal2 ;
  RECT 3445.120 500.640 3448.660 501.760 ;
  LAYER metal1 ;
  RECT 3445.120 500.640 3448.660 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3432.100 500.640 3435.640 501.760 ;
  LAYER metal4 ;
  RECT 3432.100 500.640 3435.640 501.760 ;
  LAYER metal3 ;
  RECT 3432.100 500.640 3435.640 501.760 ;
  LAYER metal2 ;
  RECT 3432.100 500.640 3435.640 501.760 ;
  LAYER metal1 ;
  RECT 3432.100 500.640 3435.640 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3418.460 500.640 3422.000 501.760 ;
  LAYER metal4 ;
  RECT 3418.460 500.640 3422.000 501.760 ;
  LAYER metal3 ;
  RECT 3418.460 500.640 3422.000 501.760 ;
  LAYER metal2 ;
  RECT 3418.460 500.640 3422.000 501.760 ;
  LAYER metal1 ;
  RECT 3418.460 500.640 3422.000 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3404.820 500.640 3408.360 501.760 ;
  LAYER metal4 ;
  RECT 3404.820 500.640 3408.360 501.760 ;
  LAYER metal3 ;
  RECT 3404.820 500.640 3408.360 501.760 ;
  LAYER metal2 ;
  RECT 3404.820 500.640 3408.360 501.760 ;
  LAYER metal1 ;
  RECT 3404.820 500.640 3408.360 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3391.800 500.640 3395.340 501.760 ;
  LAYER metal4 ;
  RECT 3391.800 500.640 3395.340 501.760 ;
  LAYER metal3 ;
  RECT 3391.800 500.640 3395.340 501.760 ;
  LAYER metal2 ;
  RECT 3391.800 500.640 3395.340 501.760 ;
  LAYER metal1 ;
  RECT 3391.800 500.640 3395.340 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3324.220 500.640 3327.760 501.760 ;
  LAYER metal4 ;
  RECT 3324.220 500.640 3327.760 501.760 ;
  LAYER metal3 ;
  RECT 3324.220 500.640 3327.760 501.760 ;
  LAYER metal2 ;
  RECT 3324.220 500.640 3327.760 501.760 ;
  LAYER metal1 ;
  RECT 3324.220 500.640 3327.760 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3311.200 500.640 3314.740 501.760 ;
  LAYER metal4 ;
  RECT 3311.200 500.640 3314.740 501.760 ;
  LAYER metal3 ;
  RECT 3311.200 500.640 3314.740 501.760 ;
  LAYER metal2 ;
  RECT 3311.200 500.640 3314.740 501.760 ;
  LAYER metal1 ;
  RECT 3311.200 500.640 3314.740 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3297.560 500.640 3301.100 501.760 ;
  LAYER metal4 ;
  RECT 3297.560 500.640 3301.100 501.760 ;
  LAYER metal3 ;
  RECT 3297.560 500.640 3301.100 501.760 ;
  LAYER metal2 ;
  RECT 3297.560 500.640 3301.100 501.760 ;
  LAYER metal1 ;
  RECT 3297.560 500.640 3301.100 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3283.920 500.640 3287.460 501.760 ;
  LAYER metal4 ;
  RECT 3283.920 500.640 3287.460 501.760 ;
  LAYER metal3 ;
  RECT 3283.920 500.640 3287.460 501.760 ;
  LAYER metal2 ;
  RECT 3283.920 500.640 3287.460 501.760 ;
  LAYER metal1 ;
  RECT 3283.920 500.640 3287.460 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3270.900 500.640 3274.440 501.760 ;
  LAYER metal4 ;
  RECT 3270.900 500.640 3274.440 501.760 ;
  LAYER metal3 ;
  RECT 3270.900 500.640 3274.440 501.760 ;
  LAYER metal2 ;
  RECT 3270.900 500.640 3274.440 501.760 ;
  LAYER metal1 ;
  RECT 3270.900 500.640 3274.440 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3257.260 500.640 3260.800 501.760 ;
  LAYER metal4 ;
  RECT 3257.260 500.640 3260.800 501.760 ;
  LAYER metal3 ;
  RECT 3257.260 500.640 3260.800 501.760 ;
  LAYER metal2 ;
  RECT 3257.260 500.640 3260.800 501.760 ;
  LAYER metal1 ;
  RECT 3257.260 500.640 3260.800 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3190.300 500.640 3193.840 501.760 ;
  LAYER metal4 ;
  RECT 3190.300 500.640 3193.840 501.760 ;
  LAYER metal3 ;
  RECT 3190.300 500.640 3193.840 501.760 ;
  LAYER metal2 ;
  RECT 3190.300 500.640 3193.840 501.760 ;
  LAYER metal1 ;
  RECT 3190.300 500.640 3193.840 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3176.660 500.640 3180.200 501.760 ;
  LAYER metal4 ;
  RECT 3176.660 500.640 3180.200 501.760 ;
  LAYER metal3 ;
  RECT 3176.660 500.640 3180.200 501.760 ;
  LAYER metal2 ;
  RECT 3176.660 500.640 3180.200 501.760 ;
  LAYER metal1 ;
  RECT 3176.660 500.640 3180.200 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3163.020 500.640 3166.560 501.760 ;
  LAYER metal4 ;
  RECT 3163.020 500.640 3166.560 501.760 ;
  LAYER metal3 ;
  RECT 3163.020 500.640 3166.560 501.760 ;
  LAYER metal2 ;
  RECT 3163.020 500.640 3166.560 501.760 ;
  LAYER metal1 ;
  RECT 3163.020 500.640 3166.560 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3149.380 500.640 3152.920 501.760 ;
  LAYER metal4 ;
  RECT 3149.380 500.640 3152.920 501.760 ;
  LAYER metal3 ;
  RECT 3149.380 500.640 3152.920 501.760 ;
  LAYER metal2 ;
  RECT 3149.380 500.640 3152.920 501.760 ;
  LAYER metal1 ;
  RECT 3149.380 500.640 3152.920 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3136.360 500.640 3139.900 501.760 ;
  LAYER metal4 ;
  RECT 3136.360 500.640 3139.900 501.760 ;
  LAYER metal3 ;
  RECT 3136.360 500.640 3139.900 501.760 ;
  LAYER metal2 ;
  RECT 3136.360 500.640 3139.900 501.760 ;
  LAYER metal1 ;
  RECT 3136.360 500.640 3139.900 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3122.720 500.640 3126.260 501.760 ;
  LAYER metal4 ;
  RECT 3122.720 500.640 3126.260 501.760 ;
  LAYER metal3 ;
  RECT 3122.720 500.640 3126.260 501.760 ;
  LAYER metal2 ;
  RECT 3122.720 500.640 3126.260 501.760 ;
  LAYER metal1 ;
  RECT 3122.720 500.640 3126.260 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3055.760 500.640 3059.300 501.760 ;
  LAYER metal4 ;
  RECT 3055.760 500.640 3059.300 501.760 ;
  LAYER metal3 ;
  RECT 3055.760 500.640 3059.300 501.760 ;
  LAYER metal2 ;
  RECT 3055.760 500.640 3059.300 501.760 ;
  LAYER metal1 ;
  RECT 3055.760 500.640 3059.300 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3042.120 500.640 3045.660 501.760 ;
  LAYER metal4 ;
  RECT 3042.120 500.640 3045.660 501.760 ;
  LAYER metal3 ;
  RECT 3042.120 500.640 3045.660 501.760 ;
  LAYER metal2 ;
  RECT 3042.120 500.640 3045.660 501.760 ;
  LAYER metal1 ;
  RECT 3042.120 500.640 3045.660 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3028.480 500.640 3032.020 501.760 ;
  LAYER metal4 ;
  RECT 3028.480 500.640 3032.020 501.760 ;
  LAYER metal3 ;
  RECT 3028.480 500.640 3032.020 501.760 ;
  LAYER metal2 ;
  RECT 3028.480 500.640 3032.020 501.760 ;
  LAYER metal1 ;
  RECT 3028.480 500.640 3032.020 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3015.460 500.640 3019.000 501.760 ;
  LAYER metal4 ;
  RECT 3015.460 500.640 3019.000 501.760 ;
  LAYER metal3 ;
  RECT 3015.460 500.640 3019.000 501.760 ;
  LAYER metal2 ;
  RECT 3015.460 500.640 3019.000 501.760 ;
  LAYER metal1 ;
  RECT 3015.460 500.640 3019.000 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3001.820 500.640 3005.360 501.760 ;
  LAYER metal4 ;
  RECT 3001.820 500.640 3005.360 501.760 ;
  LAYER metal3 ;
  RECT 3001.820 500.640 3005.360 501.760 ;
  LAYER metal2 ;
  RECT 3001.820 500.640 3005.360 501.760 ;
  LAYER metal1 ;
  RECT 3001.820 500.640 3005.360 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2988.180 500.640 2991.720 501.760 ;
  LAYER metal4 ;
  RECT 2988.180 500.640 2991.720 501.760 ;
  LAYER metal3 ;
  RECT 2988.180 500.640 2991.720 501.760 ;
  LAYER metal2 ;
  RECT 2988.180 500.640 2991.720 501.760 ;
  LAYER metal1 ;
  RECT 2988.180 500.640 2991.720 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2921.220 500.640 2924.760 501.760 ;
  LAYER metal4 ;
  RECT 2921.220 500.640 2924.760 501.760 ;
  LAYER metal3 ;
  RECT 2921.220 500.640 2924.760 501.760 ;
  LAYER metal2 ;
  RECT 2921.220 500.640 2924.760 501.760 ;
  LAYER metal1 ;
  RECT 2921.220 500.640 2924.760 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2907.580 500.640 2911.120 501.760 ;
  LAYER metal4 ;
  RECT 2907.580 500.640 2911.120 501.760 ;
  LAYER metal3 ;
  RECT 2907.580 500.640 2911.120 501.760 ;
  LAYER metal2 ;
  RECT 2907.580 500.640 2911.120 501.760 ;
  LAYER metal1 ;
  RECT 2907.580 500.640 2911.120 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2894.560 500.640 2898.100 501.760 ;
  LAYER metal4 ;
  RECT 2894.560 500.640 2898.100 501.760 ;
  LAYER metal3 ;
  RECT 2894.560 500.640 2898.100 501.760 ;
  LAYER metal2 ;
  RECT 2894.560 500.640 2898.100 501.760 ;
  LAYER metal1 ;
  RECT 2894.560 500.640 2898.100 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2880.920 500.640 2884.460 501.760 ;
  LAYER metal4 ;
  RECT 2880.920 500.640 2884.460 501.760 ;
  LAYER metal3 ;
  RECT 2880.920 500.640 2884.460 501.760 ;
  LAYER metal2 ;
  RECT 2880.920 500.640 2884.460 501.760 ;
  LAYER metal1 ;
  RECT 2880.920 500.640 2884.460 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2867.280 500.640 2870.820 501.760 ;
  LAYER metal4 ;
  RECT 2867.280 500.640 2870.820 501.760 ;
  LAYER metal3 ;
  RECT 2867.280 500.640 2870.820 501.760 ;
  LAYER metal2 ;
  RECT 2867.280 500.640 2870.820 501.760 ;
  LAYER metal1 ;
  RECT 2867.280 500.640 2870.820 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2854.260 500.640 2857.800 501.760 ;
  LAYER metal4 ;
  RECT 2854.260 500.640 2857.800 501.760 ;
  LAYER metal3 ;
  RECT 2854.260 500.640 2857.800 501.760 ;
  LAYER metal2 ;
  RECT 2854.260 500.640 2857.800 501.760 ;
  LAYER metal1 ;
  RECT 2854.260 500.640 2857.800 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2786.680 500.640 2790.220 501.760 ;
  LAYER metal4 ;
  RECT 2786.680 500.640 2790.220 501.760 ;
  LAYER metal3 ;
  RECT 2786.680 500.640 2790.220 501.760 ;
  LAYER metal2 ;
  RECT 2786.680 500.640 2790.220 501.760 ;
  LAYER metal1 ;
  RECT 2786.680 500.640 2790.220 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2773.660 500.640 2777.200 501.760 ;
  LAYER metal4 ;
  RECT 2773.660 500.640 2777.200 501.760 ;
  LAYER metal3 ;
  RECT 2773.660 500.640 2777.200 501.760 ;
  LAYER metal2 ;
  RECT 2773.660 500.640 2777.200 501.760 ;
  LAYER metal1 ;
  RECT 2773.660 500.640 2777.200 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2760.020 500.640 2763.560 501.760 ;
  LAYER metal4 ;
  RECT 2760.020 500.640 2763.560 501.760 ;
  LAYER metal3 ;
  RECT 2760.020 500.640 2763.560 501.760 ;
  LAYER metal2 ;
  RECT 2760.020 500.640 2763.560 501.760 ;
  LAYER metal1 ;
  RECT 2760.020 500.640 2763.560 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2746.380 500.640 2749.920 501.760 ;
  LAYER metal4 ;
  RECT 2746.380 500.640 2749.920 501.760 ;
  LAYER metal3 ;
  RECT 2746.380 500.640 2749.920 501.760 ;
  LAYER metal2 ;
  RECT 2746.380 500.640 2749.920 501.760 ;
  LAYER metal1 ;
  RECT 2746.380 500.640 2749.920 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2732.740 500.640 2736.280 501.760 ;
  LAYER metal4 ;
  RECT 2732.740 500.640 2736.280 501.760 ;
  LAYER metal3 ;
  RECT 2732.740 500.640 2736.280 501.760 ;
  LAYER metal2 ;
  RECT 2732.740 500.640 2736.280 501.760 ;
  LAYER metal1 ;
  RECT 2732.740 500.640 2736.280 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2719.720 500.640 2723.260 501.760 ;
  LAYER metal4 ;
  RECT 2719.720 500.640 2723.260 501.760 ;
  LAYER metal3 ;
  RECT 2719.720 500.640 2723.260 501.760 ;
  LAYER metal2 ;
  RECT 2719.720 500.640 2723.260 501.760 ;
  LAYER metal1 ;
  RECT 2719.720 500.640 2723.260 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2652.140 500.640 2655.680 501.760 ;
  LAYER metal4 ;
  RECT 2652.140 500.640 2655.680 501.760 ;
  LAYER metal3 ;
  RECT 2652.140 500.640 2655.680 501.760 ;
  LAYER metal2 ;
  RECT 2652.140 500.640 2655.680 501.760 ;
  LAYER metal1 ;
  RECT 2652.140 500.640 2655.680 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2639.120 500.640 2642.660 501.760 ;
  LAYER metal4 ;
  RECT 2639.120 500.640 2642.660 501.760 ;
  LAYER metal3 ;
  RECT 2639.120 500.640 2642.660 501.760 ;
  LAYER metal2 ;
  RECT 2639.120 500.640 2642.660 501.760 ;
  LAYER metal1 ;
  RECT 2639.120 500.640 2642.660 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2625.480 500.640 2629.020 501.760 ;
  LAYER metal4 ;
  RECT 2625.480 500.640 2629.020 501.760 ;
  LAYER metal3 ;
  RECT 2625.480 500.640 2629.020 501.760 ;
  LAYER metal2 ;
  RECT 2625.480 500.640 2629.020 501.760 ;
  LAYER metal1 ;
  RECT 2625.480 500.640 2629.020 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2611.840 500.640 2615.380 501.760 ;
  LAYER metal4 ;
  RECT 2611.840 500.640 2615.380 501.760 ;
  LAYER metal3 ;
  RECT 2611.840 500.640 2615.380 501.760 ;
  LAYER metal2 ;
  RECT 2611.840 500.640 2615.380 501.760 ;
  LAYER metal1 ;
  RECT 2611.840 500.640 2615.380 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2598.820 500.640 2602.360 501.760 ;
  LAYER metal4 ;
  RECT 2598.820 500.640 2602.360 501.760 ;
  LAYER metal3 ;
  RECT 2598.820 500.640 2602.360 501.760 ;
  LAYER metal2 ;
  RECT 2598.820 500.640 2602.360 501.760 ;
  LAYER metal1 ;
  RECT 2598.820 500.640 2602.360 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2585.180 500.640 2588.720 501.760 ;
  LAYER metal4 ;
  RECT 2585.180 500.640 2588.720 501.760 ;
  LAYER metal3 ;
  RECT 2585.180 500.640 2588.720 501.760 ;
  LAYER metal2 ;
  RECT 2585.180 500.640 2588.720 501.760 ;
  LAYER metal1 ;
  RECT 2585.180 500.640 2588.720 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2518.220 500.640 2521.760 501.760 ;
  LAYER metal4 ;
  RECT 2518.220 500.640 2521.760 501.760 ;
  LAYER metal3 ;
  RECT 2518.220 500.640 2521.760 501.760 ;
  LAYER metal2 ;
  RECT 2518.220 500.640 2521.760 501.760 ;
  LAYER metal1 ;
  RECT 2518.220 500.640 2521.760 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2504.580 500.640 2508.120 501.760 ;
  LAYER metal4 ;
  RECT 2504.580 500.640 2508.120 501.760 ;
  LAYER metal3 ;
  RECT 2504.580 500.640 2508.120 501.760 ;
  LAYER metal2 ;
  RECT 2504.580 500.640 2508.120 501.760 ;
  LAYER metal1 ;
  RECT 2504.580 500.640 2508.120 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2490.940 500.640 2494.480 501.760 ;
  LAYER metal4 ;
  RECT 2490.940 500.640 2494.480 501.760 ;
  LAYER metal3 ;
  RECT 2490.940 500.640 2494.480 501.760 ;
  LAYER metal2 ;
  RECT 2490.940 500.640 2494.480 501.760 ;
  LAYER metal1 ;
  RECT 2490.940 500.640 2494.480 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2477.920 500.640 2481.460 501.760 ;
  LAYER metal4 ;
  RECT 2477.920 500.640 2481.460 501.760 ;
  LAYER metal3 ;
  RECT 2477.920 500.640 2481.460 501.760 ;
  LAYER metal2 ;
  RECT 2477.920 500.640 2481.460 501.760 ;
  LAYER metal1 ;
  RECT 2477.920 500.640 2481.460 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2464.280 500.640 2467.820 501.760 ;
  LAYER metal4 ;
  RECT 2464.280 500.640 2467.820 501.760 ;
  LAYER metal3 ;
  RECT 2464.280 500.640 2467.820 501.760 ;
  LAYER metal2 ;
  RECT 2464.280 500.640 2467.820 501.760 ;
  LAYER metal1 ;
  RECT 2464.280 500.640 2467.820 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2450.640 500.640 2454.180 501.760 ;
  LAYER metal4 ;
  RECT 2450.640 500.640 2454.180 501.760 ;
  LAYER metal3 ;
  RECT 2450.640 500.640 2454.180 501.760 ;
  LAYER metal2 ;
  RECT 2450.640 500.640 2454.180 501.760 ;
  LAYER metal1 ;
  RECT 2450.640 500.640 2454.180 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2383.680 500.640 2387.220 501.760 ;
  LAYER metal4 ;
  RECT 2383.680 500.640 2387.220 501.760 ;
  LAYER metal3 ;
  RECT 2383.680 500.640 2387.220 501.760 ;
  LAYER metal2 ;
  RECT 2383.680 500.640 2387.220 501.760 ;
  LAYER metal1 ;
  RECT 2383.680 500.640 2387.220 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2370.040 500.640 2373.580 501.760 ;
  LAYER metal4 ;
  RECT 2370.040 500.640 2373.580 501.760 ;
  LAYER metal3 ;
  RECT 2370.040 500.640 2373.580 501.760 ;
  LAYER metal2 ;
  RECT 2370.040 500.640 2373.580 501.760 ;
  LAYER metal1 ;
  RECT 2370.040 500.640 2373.580 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2357.020 500.640 2360.560 501.760 ;
  LAYER metal4 ;
  RECT 2357.020 500.640 2360.560 501.760 ;
  LAYER metal3 ;
  RECT 2357.020 500.640 2360.560 501.760 ;
  LAYER metal2 ;
  RECT 2357.020 500.640 2360.560 501.760 ;
  LAYER metal1 ;
  RECT 2357.020 500.640 2360.560 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2343.380 500.640 2346.920 501.760 ;
  LAYER metal4 ;
  RECT 2343.380 500.640 2346.920 501.760 ;
  LAYER metal3 ;
  RECT 2343.380 500.640 2346.920 501.760 ;
  LAYER metal2 ;
  RECT 2343.380 500.640 2346.920 501.760 ;
  LAYER metal1 ;
  RECT 2343.380 500.640 2346.920 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2329.740 500.640 2333.280 501.760 ;
  LAYER metal4 ;
  RECT 2329.740 500.640 2333.280 501.760 ;
  LAYER metal3 ;
  RECT 2329.740 500.640 2333.280 501.760 ;
  LAYER metal2 ;
  RECT 2329.740 500.640 2333.280 501.760 ;
  LAYER metal1 ;
  RECT 2329.740 500.640 2333.280 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2316.100 500.640 2319.640 501.760 ;
  LAYER metal4 ;
  RECT 2316.100 500.640 2319.640 501.760 ;
  LAYER metal3 ;
  RECT 2316.100 500.640 2319.640 501.760 ;
  LAYER metal2 ;
  RECT 2316.100 500.640 2319.640 501.760 ;
  LAYER metal1 ;
  RECT 2316.100 500.640 2319.640 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2249.140 500.640 2252.680 501.760 ;
  LAYER metal4 ;
  RECT 2249.140 500.640 2252.680 501.760 ;
  LAYER metal3 ;
  RECT 2249.140 500.640 2252.680 501.760 ;
  LAYER metal2 ;
  RECT 2249.140 500.640 2252.680 501.760 ;
  LAYER metal1 ;
  RECT 2249.140 500.640 2252.680 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2235.500 500.640 2239.040 501.760 ;
  LAYER metal4 ;
  RECT 2235.500 500.640 2239.040 501.760 ;
  LAYER metal3 ;
  RECT 2235.500 500.640 2239.040 501.760 ;
  LAYER metal2 ;
  RECT 2235.500 500.640 2239.040 501.760 ;
  LAYER metal1 ;
  RECT 2235.500 500.640 2239.040 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2222.480 500.640 2226.020 501.760 ;
  LAYER metal4 ;
  RECT 2222.480 500.640 2226.020 501.760 ;
  LAYER metal3 ;
  RECT 2222.480 500.640 2226.020 501.760 ;
  LAYER metal2 ;
  RECT 2222.480 500.640 2226.020 501.760 ;
  LAYER metal1 ;
  RECT 2222.480 500.640 2226.020 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2208.840 500.640 2212.380 501.760 ;
  LAYER metal4 ;
  RECT 2208.840 500.640 2212.380 501.760 ;
  LAYER metal3 ;
  RECT 2208.840 500.640 2212.380 501.760 ;
  LAYER metal2 ;
  RECT 2208.840 500.640 2212.380 501.760 ;
  LAYER metal1 ;
  RECT 2208.840 500.640 2212.380 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2195.200 500.640 2198.740 501.760 ;
  LAYER metal4 ;
  RECT 2195.200 500.640 2198.740 501.760 ;
  LAYER metal3 ;
  RECT 2195.200 500.640 2198.740 501.760 ;
  LAYER metal2 ;
  RECT 2195.200 500.640 2198.740 501.760 ;
  LAYER metal1 ;
  RECT 2195.200 500.640 2198.740 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2182.180 500.640 2185.720 501.760 ;
  LAYER metal4 ;
  RECT 2182.180 500.640 2185.720 501.760 ;
  LAYER metal3 ;
  RECT 2182.180 500.640 2185.720 501.760 ;
  LAYER metal2 ;
  RECT 2182.180 500.640 2185.720 501.760 ;
  LAYER metal1 ;
  RECT 2182.180 500.640 2185.720 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2114.600 500.640 2118.140 501.760 ;
  LAYER metal4 ;
  RECT 2114.600 500.640 2118.140 501.760 ;
  LAYER metal3 ;
  RECT 2114.600 500.640 2118.140 501.760 ;
  LAYER metal2 ;
  RECT 2114.600 500.640 2118.140 501.760 ;
  LAYER metal1 ;
  RECT 2114.600 500.640 2118.140 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2101.580 500.640 2105.120 501.760 ;
  LAYER metal4 ;
  RECT 2101.580 500.640 2105.120 501.760 ;
  LAYER metal3 ;
  RECT 2101.580 500.640 2105.120 501.760 ;
  LAYER metal2 ;
  RECT 2101.580 500.640 2105.120 501.760 ;
  LAYER metal1 ;
  RECT 2101.580 500.640 2105.120 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2087.940 500.640 2091.480 501.760 ;
  LAYER metal4 ;
  RECT 2087.940 500.640 2091.480 501.760 ;
  LAYER metal3 ;
  RECT 2087.940 500.640 2091.480 501.760 ;
  LAYER metal2 ;
  RECT 2087.940 500.640 2091.480 501.760 ;
  LAYER metal1 ;
  RECT 2087.940 500.640 2091.480 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2074.300 500.640 2077.840 501.760 ;
  LAYER metal4 ;
  RECT 2074.300 500.640 2077.840 501.760 ;
  LAYER metal3 ;
  RECT 2074.300 500.640 2077.840 501.760 ;
  LAYER metal2 ;
  RECT 2074.300 500.640 2077.840 501.760 ;
  LAYER metal1 ;
  RECT 2074.300 500.640 2077.840 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2061.280 500.640 2064.820 501.760 ;
  LAYER metal4 ;
  RECT 2061.280 500.640 2064.820 501.760 ;
  LAYER metal3 ;
  RECT 2061.280 500.640 2064.820 501.760 ;
  LAYER metal2 ;
  RECT 2061.280 500.640 2064.820 501.760 ;
  LAYER metal1 ;
  RECT 2061.280 500.640 2064.820 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2047.640 500.640 2051.180 501.760 ;
  LAYER metal4 ;
  RECT 2047.640 500.640 2051.180 501.760 ;
  LAYER metal3 ;
  RECT 2047.640 500.640 2051.180 501.760 ;
  LAYER metal2 ;
  RECT 2047.640 500.640 2051.180 501.760 ;
  LAYER metal1 ;
  RECT 2047.640 500.640 2051.180 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1980.680 500.640 1984.220 501.760 ;
  LAYER metal4 ;
  RECT 1980.680 500.640 1984.220 501.760 ;
  LAYER metal3 ;
  RECT 1980.680 500.640 1984.220 501.760 ;
  LAYER metal2 ;
  RECT 1980.680 500.640 1984.220 501.760 ;
  LAYER metal1 ;
  RECT 1980.680 500.640 1984.220 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1967.040 500.640 1970.580 501.760 ;
  LAYER metal4 ;
  RECT 1967.040 500.640 1970.580 501.760 ;
  LAYER metal3 ;
  RECT 1967.040 500.640 1970.580 501.760 ;
  LAYER metal2 ;
  RECT 1967.040 500.640 1970.580 501.760 ;
  LAYER metal1 ;
  RECT 1967.040 500.640 1970.580 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1953.400 500.640 1956.940 501.760 ;
  LAYER metal4 ;
  RECT 1953.400 500.640 1956.940 501.760 ;
  LAYER metal3 ;
  RECT 1953.400 500.640 1956.940 501.760 ;
  LAYER metal2 ;
  RECT 1953.400 500.640 1956.940 501.760 ;
  LAYER metal1 ;
  RECT 1953.400 500.640 1956.940 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1940.380 500.640 1943.920 501.760 ;
  LAYER metal4 ;
  RECT 1940.380 500.640 1943.920 501.760 ;
  LAYER metal3 ;
  RECT 1940.380 500.640 1943.920 501.760 ;
  LAYER metal2 ;
  RECT 1940.380 500.640 1943.920 501.760 ;
  LAYER metal1 ;
  RECT 1940.380 500.640 1943.920 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1926.740 500.640 1930.280 501.760 ;
  LAYER metal4 ;
  RECT 1926.740 500.640 1930.280 501.760 ;
  LAYER metal3 ;
  RECT 1926.740 500.640 1930.280 501.760 ;
  LAYER metal2 ;
  RECT 1926.740 500.640 1930.280 501.760 ;
  LAYER metal1 ;
  RECT 1926.740 500.640 1930.280 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1913.100 500.640 1916.640 501.760 ;
  LAYER metal4 ;
  RECT 1913.100 500.640 1916.640 501.760 ;
  LAYER metal3 ;
  RECT 1913.100 500.640 1916.640 501.760 ;
  LAYER metal2 ;
  RECT 1913.100 500.640 1916.640 501.760 ;
  LAYER metal1 ;
  RECT 1913.100 500.640 1916.640 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1850.480 500.640 1854.020 501.760 ;
  LAYER metal4 ;
  RECT 1850.480 500.640 1854.020 501.760 ;
  LAYER metal3 ;
  RECT 1850.480 500.640 1854.020 501.760 ;
  LAYER metal2 ;
  RECT 1850.480 500.640 1854.020 501.760 ;
  LAYER metal1 ;
  RECT 1850.480 500.640 1854.020 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1841.800 500.640 1845.340 501.760 ;
  LAYER metal4 ;
  RECT 1841.800 500.640 1845.340 501.760 ;
  LAYER metal3 ;
  RECT 1841.800 500.640 1845.340 501.760 ;
  LAYER metal2 ;
  RECT 1841.800 500.640 1845.340 501.760 ;
  LAYER metal1 ;
  RECT 1841.800 500.640 1845.340 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1828.780 500.640 1832.320 501.760 ;
  LAYER metal4 ;
  RECT 1828.780 500.640 1832.320 501.760 ;
  LAYER metal3 ;
  RECT 1828.780 500.640 1832.320 501.760 ;
  LAYER metal2 ;
  RECT 1828.780 500.640 1832.320 501.760 ;
  LAYER metal1 ;
  RECT 1828.780 500.640 1832.320 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1784.140 500.640 1787.680 501.760 ;
  LAYER metal4 ;
  RECT 1784.140 500.640 1787.680 501.760 ;
  LAYER metal3 ;
  RECT 1784.140 500.640 1787.680 501.760 ;
  LAYER metal2 ;
  RECT 1784.140 500.640 1787.680 501.760 ;
  LAYER metal1 ;
  RECT 1784.140 500.640 1787.680 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1761.200 500.640 1764.740 501.760 ;
  LAYER metal4 ;
  RECT 1761.200 500.640 1764.740 501.760 ;
  LAYER metal3 ;
  RECT 1761.200 500.640 1764.740 501.760 ;
  LAYER metal2 ;
  RECT 1761.200 500.640 1764.740 501.760 ;
  LAYER metal1 ;
  RECT 1761.200 500.640 1764.740 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1752.520 500.640 1756.060 501.760 ;
  LAYER metal4 ;
  RECT 1752.520 500.640 1756.060 501.760 ;
  LAYER metal3 ;
  RECT 1752.520 500.640 1756.060 501.760 ;
  LAYER metal2 ;
  RECT 1752.520 500.640 1756.060 501.760 ;
  LAYER metal1 ;
  RECT 1752.520 500.640 1756.060 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1694.860 500.640 1698.400 501.760 ;
  LAYER metal4 ;
  RECT 1694.860 500.640 1698.400 501.760 ;
  LAYER metal3 ;
  RECT 1694.860 500.640 1698.400 501.760 ;
  LAYER metal2 ;
  RECT 1694.860 500.640 1698.400 501.760 ;
  LAYER metal1 ;
  RECT 1694.860 500.640 1698.400 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1681.220 500.640 1684.760 501.760 ;
  LAYER metal4 ;
  RECT 1681.220 500.640 1684.760 501.760 ;
  LAYER metal3 ;
  RECT 1681.220 500.640 1684.760 501.760 ;
  LAYER metal2 ;
  RECT 1681.220 500.640 1684.760 501.760 ;
  LAYER metal1 ;
  RECT 1681.220 500.640 1684.760 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1668.200 500.640 1671.740 501.760 ;
  LAYER metal4 ;
  RECT 1668.200 500.640 1671.740 501.760 ;
  LAYER metal3 ;
  RECT 1668.200 500.640 1671.740 501.760 ;
  LAYER metal2 ;
  RECT 1668.200 500.640 1671.740 501.760 ;
  LAYER metal1 ;
  RECT 1668.200 500.640 1671.740 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1654.560 500.640 1658.100 501.760 ;
  LAYER metal4 ;
  RECT 1654.560 500.640 1658.100 501.760 ;
  LAYER metal3 ;
  RECT 1654.560 500.640 1658.100 501.760 ;
  LAYER metal2 ;
  RECT 1654.560 500.640 1658.100 501.760 ;
  LAYER metal1 ;
  RECT 1654.560 500.640 1658.100 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1640.920 500.640 1644.460 501.760 ;
  LAYER metal4 ;
  RECT 1640.920 500.640 1644.460 501.760 ;
  LAYER metal3 ;
  RECT 1640.920 500.640 1644.460 501.760 ;
  LAYER metal2 ;
  RECT 1640.920 500.640 1644.460 501.760 ;
  LAYER metal1 ;
  RECT 1640.920 500.640 1644.460 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1627.900 500.640 1631.440 501.760 ;
  LAYER metal4 ;
  RECT 1627.900 500.640 1631.440 501.760 ;
  LAYER metal3 ;
  RECT 1627.900 500.640 1631.440 501.760 ;
  LAYER metal2 ;
  RECT 1627.900 500.640 1631.440 501.760 ;
  LAYER metal1 ;
  RECT 1627.900 500.640 1631.440 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1560.320 500.640 1563.860 501.760 ;
  LAYER metal4 ;
  RECT 1560.320 500.640 1563.860 501.760 ;
  LAYER metal3 ;
  RECT 1560.320 500.640 1563.860 501.760 ;
  LAYER metal2 ;
  RECT 1560.320 500.640 1563.860 501.760 ;
  LAYER metal1 ;
  RECT 1560.320 500.640 1563.860 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1547.300 500.640 1550.840 501.760 ;
  LAYER metal4 ;
  RECT 1547.300 500.640 1550.840 501.760 ;
  LAYER metal3 ;
  RECT 1547.300 500.640 1550.840 501.760 ;
  LAYER metal2 ;
  RECT 1547.300 500.640 1550.840 501.760 ;
  LAYER metal1 ;
  RECT 1547.300 500.640 1550.840 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1533.660 500.640 1537.200 501.760 ;
  LAYER metal4 ;
  RECT 1533.660 500.640 1537.200 501.760 ;
  LAYER metal3 ;
  RECT 1533.660 500.640 1537.200 501.760 ;
  LAYER metal2 ;
  RECT 1533.660 500.640 1537.200 501.760 ;
  LAYER metal1 ;
  RECT 1533.660 500.640 1537.200 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1520.020 500.640 1523.560 501.760 ;
  LAYER metal4 ;
  RECT 1520.020 500.640 1523.560 501.760 ;
  LAYER metal3 ;
  RECT 1520.020 500.640 1523.560 501.760 ;
  LAYER metal2 ;
  RECT 1520.020 500.640 1523.560 501.760 ;
  LAYER metal1 ;
  RECT 1520.020 500.640 1523.560 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1507.000 500.640 1510.540 501.760 ;
  LAYER metal4 ;
  RECT 1507.000 500.640 1510.540 501.760 ;
  LAYER metal3 ;
  RECT 1507.000 500.640 1510.540 501.760 ;
  LAYER metal2 ;
  RECT 1507.000 500.640 1510.540 501.760 ;
  LAYER metal1 ;
  RECT 1507.000 500.640 1510.540 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1493.360 500.640 1496.900 501.760 ;
  LAYER metal4 ;
  RECT 1493.360 500.640 1496.900 501.760 ;
  LAYER metal3 ;
  RECT 1493.360 500.640 1496.900 501.760 ;
  LAYER metal2 ;
  RECT 1493.360 500.640 1496.900 501.760 ;
  LAYER metal1 ;
  RECT 1493.360 500.640 1496.900 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1426.400 500.640 1429.940 501.760 ;
  LAYER metal4 ;
  RECT 1426.400 500.640 1429.940 501.760 ;
  LAYER metal3 ;
  RECT 1426.400 500.640 1429.940 501.760 ;
  LAYER metal2 ;
  RECT 1426.400 500.640 1429.940 501.760 ;
  LAYER metal1 ;
  RECT 1426.400 500.640 1429.940 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1412.760 500.640 1416.300 501.760 ;
  LAYER metal4 ;
  RECT 1412.760 500.640 1416.300 501.760 ;
  LAYER metal3 ;
  RECT 1412.760 500.640 1416.300 501.760 ;
  LAYER metal2 ;
  RECT 1412.760 500.640 1416.300 501.760 ;
  LAYER metal1 ;
  RECT 1412.760 500.640 1416.300 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1399.120 500.640 1402.660 501.760 ;
  LAYER metal4 ;
  RECT 1399.120 500.640 1402.660 501.760 ;
  LAYER metal3 ;
  RECT 1399.120 500.640 1402.660 501.760 ;
  LAYER metal2 ;
  RECT 1399.120 500.640 1402.660 501.760 ;
  LAYER metal1 ;
  RECT 1399.120 500.640 1402.660 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1386.100 500.640 1389.640 501.760 ;
  LAYER metal4 ;
  RECT 1386.100 500.640 1389.640 501.760 ;
  LAYER metal3 ;
  RECT 1386.100 500.640 1389.640 501.760 ;
  LAYER metal2 ;
  RECT 1386.100 500.640 1389.640 501.760 ;
  LAYER metal1 ;
  RECT 1386.100 500.640 1389.640 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1372.460 500.640 1376.000 501.760 ;
  LAYER metal4 ;
  RECT 1372.460 500.640 1376.000 501.760 ;
  LAYER metal3 ;
  RECT 1372.460 500.640 1376.000 501.760 ;
  LAYER metal2 ;
  RECT 1372.460 500.640 1376.000 501.760 ;
  LAYER metal1 ;
  RECT 1372.460 500.640 1376.000 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1358.820 500.640 1362.360 501.760 ;
  LAYER metal4 ;
  RECT 1358.820 500.640 1362.360 501.760 ;
  LAYER metal3 ;
  RECT 1358.820 500.640 1362.360 501.760 ;
  LAYER metal2 ;
  RECT 1358.820 500.640 1362.360 501.760 ;
  LAYER metal1 ;
  RECT 1358.820 500.640 1362.360 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1291.860 500.640 1295.400 501.760 ;
  LAYER metal4 ;
  RECT 1291.860 500.640 1295.400 501.760 ;
  LAYER metal3 ;
  RECT 1291.860 500.640 1295.400 501.760 ;
  LAYER metal2 ;
  RECT 1291.860 500.640 1295.400 501.760 ;
  LAYER metal1 ;
  RECT 1291.860 500.640 1295.400 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1278.220 500.640 1281.760 501.760 ;
  LAYER metal4 ;
  RECT 1278.220 500.640 1281.760 501.760 ;
  LAYER metal3 ;
  RECT 1278.220 500.640 1281.760 501.760 ;
  LAYER metal2 ;
  RECT 1278.220 500.640 1281.760 501.760 ;
  LAYER metal1 ;
  RECT 1278.220 500.640 1281.760 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1264.580 500.640 1268.120 501.760 ;
  LAYER metal4 ;
  RECT 1264.580 500.640 1268.120 501.760 ;
  LAYER metal3 ;
  RECT 1264.580 500.640 1268.120 501.760 ;
  LAYER metal2 ;
  RECT 1264.580 500.640 1268.120 501.760 ;
  LAYER metal1 ;
  RECT 1264.580 500.640 1268.120 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1251.560 500.640 1255.100 501.760 ;
  LAYER metal4 ;
  RECT 1251.560 500.640 1255.100 501.760 ;
  LAYER metal3 ;
  RECT 1251.560 500.640 1255.100 501.760 ;
  LAYER metal2 ;
  RECT 1251.560 500.640 1255.100 501.760 ;
  LAYER metal1 ;
  RECT 1251.560 500.640 1255.100 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1237.920 500.640 1241.460 501.760 ;
  LAYER metal4 ;
  RECT 1237.920 500.640 1241.460 501.760 ;
  LAYER metal3 ;
  RECT 1237.920 500.640 1241.460 501.760 ;
  LAYER metal2 ;
  RECT 1237.920 500.640 1241.460 501.760 ;
  LAYER metal1 ;
  RECT 1237.920 500.640 1241.460 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1224.280 500.640 1227.820 501.760 ;
  LAYER metal4 ;
  RECT 1224.280 500.640 1227.820 501.760 ;
  LAYER metal3 ;
  RECT 1224.280 500.640 1227.820 501.760 ;
  LAYER metal2 ;
  RECT 1224.280 500.640 1227.820 501.760 ;
  LAYER metal1 ;
  RECT 1224.280 500.640 1227.820 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1157.320 500.640 1160.860 501.760 ;
  LAYER metal4 ;
  RECT 1157.320 500.640 1160.860 501.760 ;
  LAYER metal3 ;
  RECT 1157.320 500.640 1160.860 501.760 ;
  LAYER metal2 ;
  RECT 1157.320 500.640 1160.860 501.760 ;
  LAYER metal1 ;
  RECT 1157.320 500.640 1160.860 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1143.680 500.640 1147.220 501.760 ;
  LAYER metal4 ;
  RECT 1143.680 500.640 1147.220 501.760 ;
  LAYER metal3 ;
  RECT 1143.680 500.640 1147.220 501.760 ;
  LAYER metal2 ;
  RECT 1143.680 500.640 1147.220 501.760 ;
  LAYER metal1 ;
  RECT 1143.680 500.640 1147.220 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1130.660 500.640 1134.200 501.760 ;
  LAYER metal4 ;
  RECT 1130.660 500.640 1134.200 501.760 ;
  LAYER metal3 ;
  RECT 1130.660 500.640 1134.200 501.760 ;
  LAYER metal2 ;
  RECT 1130.660 500.640 1134.200 501.760 ;
  LAYER metal1 ;
  RECT 1130.660 500.640 1134.200 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1117.020 500.640 1120.560 501.760 ;
  LAYER metal4 ;
  RECT 1117.020 500.640 1120.560 501.760 ;
  LAYER metal3 ;
  RECT 1117.020 500.640 1120.560 501.760 ;
  LAYER metal2 ;
  RECT 1117.020 500.640 1120.560 501.760 ;
  LAYER metal1 ;
  RECT 1117.020 500.640 1120.560 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1103.380 500.640 1106.920 501.760 ;
  LAYER metal4 ;
  RECT 1103.380 500.640 1106.920 501.760 ;
  LAYER metal3 ;
  RECT 1103.380 500.640 1106.920 501.760 ;
  LAYER metal2 ;
  RECT 1103.380 500.640 1106.920 501.760 ;
  LAYER metal1 ;
  RECT 1103.380 500.640 1106.920 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1090.360 500.640 1093.900 501.760 ;
  LAYER metal4 ;
  RECT 1090.360 500.640 1093.900 501.760 ;
  LAYER metal3 ;
  RECT 1090.360 500.640 1093.900 501.760 ;
  LAYER metal2 ;
  RECT 1090.360 500.640 1093.900 501.760 ;
  LAYER metal1 ;
  RECT 1090.360 500.640 1093.900 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1022.780 500.640 1026.320 501.760 ;
  LAYER metal4 ;
  RECT 1022.780 500.640 1026.320 501.760 ;
  LAYER metal3 ;
  RECT 1022.780 500.640 1026.320 501.760 ;
  LAYER metal2 ;
  RECT 1022.780 500.640 1026.320 501.760 ;
  LAYER metal1 ;
  RECT 1022.780 500.640 1026.320 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1009.760 500.640 1013.300 501.760 ;
  LAYER metal4 ;
  RECT 1009.760 500.640 1013.300 501.760 ;
  LAYER metal3 ;
  RECT 1009.760 500.640 1013.300 501.760 ;
  LAYER metal2 ;
  RECT 1009.760 500.640 1013.300 501.760 ;
  LAYER metal1 ;
  RECT 1009.760 500.640 1013.300 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 996.120 500.640 999.660 501.760 ;
  LAYER metal4 ;
  RECT 996.120 500.640 999.660 501.760 ;
  LAYER metal3 ;
  RECT 996.120 500.640 999.660 501.760 ;
  LAYER metal2 ;
  RECT 996.120 500.640 999.660 501.760 ;
  LAYER metal1 ;
  RECT 996.120 500.640 999.660 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 982.480 500.640 986.020 501.760 ;
  LAYER metal4 ;
  RECT 982.480 500.640 986.020 501.760 ;
  LAYER metal3 ;
  RECT 982.480 500.640 986.020 501.760 ;
  LAYER metal2 ;
  RECT 982.480 500.640 986.020 501.760 ;
  LAYER metal1 ;
  RECT 982.480 500.640 986.020 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 969.460 500.640 973.000 501.760 ;
  LAYER metal4 ;
  RECT 969.460 500.640 973.000 501.760 ;
  LAYER metal3 ;
  RECT 969.460 500.640 973.000 501.760 ;
  LAYER metal2 ;
  RECT 969.460 500.640 973.000 501.760 ;
  LAYER metal1 ;
  RECT 969.460 500.640 973.000 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 955.820 500.640 959.360 501.760 ;
  LAYER metal4 ;
  RECT 955.820 500.640 959.360 501.760 ;
  LAYER metal3 ;
  RECT 955.820 500.640 959.360 501.760 ;
  LAYER metal2 ;
  RECT 955.820 500.640 959.360 501.760 ;
  LAYER metal1 ;
  RECT 955.820 500.640 959.360 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 888.240 500.640 891.780 501.760 ;
  LAYER metal4 ;
  RECT 888.240 500.640 891.780 501.760 ;
  LAYER metal3 ;
  RECT 888.240 500.640 891.780 501.760 ;
  LAYER metal2 ;
  RECT 888.240 500.640 891.780 501.760 ;
  LAYER metal1 ;
  RECT 888.240 500.640 891.780 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 875.220 500.640 878.760 501.760 ;
  LAYER metal4 ;
  RECT 875.220 500.640 878.760 501.760 ;
  LAYER metal3 ;
  RECT 875.220 500.640 878.760 501.760 ;
  LAYER metal2 ;
  RECT 875.220 500.640 878.760 501.760 ;
  LAYER metal1 ;
  RECT 875.220 500.640 878.760 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 861.580 500.640 865.120 501.760 ;
  LAYER metal4 ;
  RECT 861.580 500.640 865.120 501.760 ;
  LAYER metal3 ;
  RECT 861.580 500.640 865.120 501.760 ;
  LAYER metal2 ;
  RECT 861.580 500.640 865.120 501.760 ;
  LAYER metal1 ;
  RECT 861.580 500.640 865.120 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 847.940 500.640 851.480 501.760 ;
  LAYER metal4 ;
  RECT 847.940 500.640 851.480 501.760 ;
  LAYER metal3 ;
  RECT 847.940 500.640 851.480 501.760 ;
  LAYER metal2 ;
  RECT 847.940 500.640 851.480 501.760 ;
  LAYER metal1 ;
  RECT 847.940 500.640 851.480 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 834.920 500.640 838.460 501.760 ;
  LAYER metal4 ;
  RECT 834.920 500.640 838.460 501.760 ;
  LAYER metal3 ;
  RECT 834.920 500.640 838.460 501.760 ;
  LAYER metal2 ;
  RECT 834.920 500.640 838.460 501.760 ;
  LAYER metal1 ;
  RECT 834.920 500.640 838.460 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 821.280 500.640 824.820 501.760 ;
  LAYER metal4 ;
  RECT 821.280 500.640 824.820 501.760 ;
  LAYER metal3 ;
  RECT 821.280 500.640 824.820 501.760 ;
  LAYER metal2 ;
  RECT 821.280 500.640 824.820 501.760 ;
  LAYER metal1 ;
  RECT 821.280 500.640 824.820 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 754.320 500.640 757.860 501.760 ;
  LAYER metal4 ;
  RECT 754.320 500.640 757.860 501.760 ;
  LAYER metal3 ;
  RECT 754.320 500.640 757.860 501.760 ;
  LAYER metal2 ;
  RECT 754.320 500.640 757.860 501.760 ;
  LAYER metal1 ;
  RECT 754.320 500.640 757.860 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 740.680 500.640 744.220 501.760 ;
  LAYER metal4 ;
  RECT 740.680 500.640 744.220 501.760 ;
  LAYER metal3 ;
  RECT 740.680 500.640 744.220 501.760 ;
  LAYER metal2 ;
  RECT 740.680 500.640 744.220 501.760 ;
  LAYER metal1 ;
  RECT 740.680 500.640 744.220 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 727.040 500.640 730.580 501.760 ;
  LAYER metal4 ;
  RECT 727.040 500.640 730.580 501.760 ;
  LAYER metal3 ;
  RECT 727.040 500.640 730.580 501.760 ;
  LAYER metal2 ;
  RECT 727.040 500.640 730.580 501.760 ;
  LAYER metal1 ;
  RECT 727.040 500.640 730.580 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 714.020 500.640 717.560 501.760 ;
  LAYER metal4 ;
  RECT 714.020 500.640 717.560 501.760 ;
  LAYER metal3 ;
  RECT 714.020 500.640 717.560 501.760 ;
  LAYER metal2 ;
  RECT 714.020 500.640 717.560 501.760 ;
  LAYER metal1 ;
  RECT 714.020 500.640 717.560 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 700.380 500.640 703.920 501.760 ;
  LAYER metal4 ;
  RECT 700.380 500.640 703.920 501.760 ;
  LAYER metal3 ;
  RECT 700.380 500.640 703.920 501.760 ;
  LAYER metal2 ;
  RECT 700.380 500.640 703.920 501.760 ;
  LAYER metal1 ;
  RECT 700.380 500.640 703.920 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 686.740 500.640 690.280 501.760 ;
  LAYER metal4 ;
  RECT 686.740 500.640 690.280 501.760 ;
  LAYER metal3 ;
  RECT 686.740 500.640 690.280 501.760 ;
  LAYER metal2 ;
  RECT 686.740 500.640 690.280 501.760 ;
  LAYER metal1 ;
  RECT 686.740 500.640 690.280 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 619.780 500.640 623.320 501.760 ;
  LAYER metal4 ;
  RECT 619.780 500.640 623.320 501.760 ;
  LAYER metal3 ;
  RECT 619.780 500.640 623.320 501.760 ;
  LAYER metal2 ;
  RECT 619.780 500.640 623.320 501.760 ;
  LAYER metal1 ;
  RECT 619.780 500.640 623.320 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 606.140 500.640 609.680 501.760 ;
  LAYER metal4 ;
  RECT 606.140 500.640 609.680 501.760 ;
  LAYER metal3 ;
  RECT 606.140 500.640 609.680 501.760 ;
  LAYER metal2 ;
  RECT 606.140 500.640 609.680 501.760 ;
  LAYER metal1 ;
  RECT 606.140 500.640 609.680 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 593.120 500.640 596.660 501.760 ;
  LAYER metal4 ;
  RECT 593.120 500.640 596.660 501.760 ;
  LAYER metal3 ;
  RECT 593.120 500.640 596.660 501.760 ;
  LAYER metal2 ;
  RECT 593.120 500.640 596.660 501.760 ;
  LAYER metal1 ;
  RECT 593.120 500.640 596.660 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 579.480 500.640 583.020 501.760 ;
  LAYER metal4 ;
  RECT 579.480 500.640 583.020 501.760 ;
  LAYER metal3 ;
  RECT 579.480 500.640 583.020 501.760 ;
  LAYER metal2 ;
  RECT 579.480 500.640 583.020 501.760 ;
  LAYER metal1 ;
  RECT 579.480 500.640 583.020 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 565.840 500.640 569.380 501.760 ;
  LAYER metal4 ;
  RECT 565.840 500.640 569.380 501.760 ;
  LAYER metal3 ;
  RECT 565.840 500.640 569.380 501.760 ;
  LAYER metal2 ;
  RECT 565.840 500.640 569.380 501.760 ;
  LAYER metal1 ;
  RECT 565.840 500.640 569.380 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 552.820 500.640 556.360 501.760 ;
  LAYER metal4 ;
  RECT 552.820 500.640 556.360 501.760 ;
  LAYER metal3 ;
  RECT 552.820 500.640 556.360 501.760 ;
  LAYER metal2 ;
  RECT 552.820 500.640 556.360 501.760 ;
  LAYER metal1 ;
  RECT 552.820 500.640 556.360 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 485.240 500.640 488.780 501.760 ;
  LAYER metal4 ;
  RECT 485.240 500.640 488.780 501.760 ;
  LAYER metal3 ;
  RECT 485.240 500.640 488.780 501.760 ;
  LAYER metal2 ;
  RECT 485.240 500.640 488.780 501.760 ;
  LAYER metal1 ;
  RECT 485.240 500.640 488.780 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 471.600 500.640 475.140 501.760 ;
  LAYER metal4 ;
  RECT 471.600 500.640 475.140 501.760 ;
  LAYER metal3 ;
  RECT 471.600 500.640 475.140 501.760 ;
  LAYER metal2 ;
  RECT 471.600 500.640 475.140 501.760 ;
  LAYER metal1 ;
  RECT 471.600 500.640 475.140 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 458.580 500.640 462.120 501.760 ;
  LAYER metal4 ;
  RECT 458.580 500.640 462.120 501.760 ;
  LAYER metal3 ;
  RECT 458.580 500.640 462.120 501.760 ;
  LAYER metal2 ;
  RECT 458.580 500.640 462.120 501.760 ;
  LAYER metal1 ;
  RECT 458.580 500.640 462.120 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 444.940 500.640 448.480 501.760 ;
  LAYER metal4 ;
  RECT 444.940 500.640 448.480 501.760 ;
  LAYER metal3 ;
  RECT 444.940 500.640 448.480 501.760 ;
  LAYER metal2 ;
  RECT 444.940 500.640 448.480 501.760 ;
  LAYER metal1 ;
  RECT 444.940 500.640 448.480 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 431.300 500.640 434.840 501.760 ;
  LAYER metal4 ;
  RECT 431.300 500.640 434.840 501.760 ;
  LAYER metal3 ;
  RECT 431.300 500.640 434.840 501.760 ;
  LAYER metal2 ;
  RECT 431.300 500.640 434.840 501.760 ;
  LAYER metal1 ;
  RECT 431.300 500.640 434.840 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 418.280 500.640 421.820 501.760 ;
  LAYER metal4 ;
  RECT 418.280 500.640 421.820 501.760 ;
  LAYER metal3 ;
  RECT 418.280 500.640 421.820 501.760 ;
  LAYER metal2 ;
  RECT 418.280 500.640 421.820 501.760 ;
  LAYER metal1 ;
  RECT 418.280 500.640 421.820 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 350.700 500.640 354.240 501.760 ;
  LAYER metal4 ;
  RECT 350.700 500.640 354.240 501.760 ;
  LAYER metal3 ;
  RECT 350.700 500.640 354.240 501.760 ;
  LAYER metal2 ;
  RECT 350.700 500.640 354.240 501.760 ;
  LAYER metal1 ;
  RECT 350.700 500.640 354.240 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 337.680 500.640 341.220 501.760 ;
  LAYER metal4 ;
  RECT 337.680 500.640 341.220 501.760 ;
  LAYER metal3 ;
  RECT 337.680 500.640 341.220 501.760 ;
  LAYER metal2 ;
  RECT 337.680 500.640 341.220 501.760 ;
  LAYER metal1 ;
  RECT 337.680 500.640 341.220 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 324.040 500.640 327.580 501.760 ;
  LAYER metal4 ;
  RECT 324.040 500.640 327.580 501.760 ;
  LAYER metal3 ;
  RECT 324.040 500.640 327.580 501.760 ;
  LAYER metal2 ;
  RECT 324.040 500.640 327.580 501.760 ;
  LAYER metal1 ;
  RECT 324.040 500.640 327.580 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 310.400 500.640 313.940 501.760 ;
  LAYER metal4 ;
  RECT 310.400 500.640 313.940 501.760 ;
  LAYER metal3 ;
  RECT 310.400 500.640 313.940 501.760 ;
  LAYER metal2 ;
  RECT 310.400 500.640 313.940 501.760 ;
  LAYER metal1 ;
  RECT 310.400 500.640 313.940 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 297.380 500.640 300.920 501.760 ;
  LAYER metal4 ;
  RECT 297.380 500.640 300.920 501.760 ;
  LAYER metal3 ;
  RECT 297.380 500.640 300.920 501.760 ;
  LAYER metal2 ;
  RECT 297.380 500.640 300.920 501.760 ;
  LAYER metal1 ;
  RECT 297.380 500.640 300.920 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 283.740 500.640 287.280 501.760 ;
  LAYER metal4 ;
  RECT 283.740 500.640 287.280 501.760 ;
  LAYER metal3 ;
  RECT 283.740 500.640 287.280 501.760 ;
  LAYER metal2 ;
  RECT 283.740 500.640 287.280 501.760 ;
  LAYER metal1 ;
  RECT 283.740 500.640 287.280 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 216.780 500.640 220.320 501.760 ;
  LAYER metal4 ;
  RECT 216.780 500.640 220.320 501.760 ;
  LAYER metal3 ;
  RECT 216.780 500.640 220.320 501.760 ;
  LAYER metal2 ;
  RECT 216.780 500.640 220.320 501.760 ;
  LAYER metal1 ;
  RECT 216.780 500.640 220.320 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 203.140 500.640 206.680 501.760 ;
  LAYER metal4 ;
  RECT 203.140 500.640 206.680 501.760 ;
  LAYER metal3 ;
  RECT 203.140 500.640 206.680 501.760 ;
  LAYER metal2 ;
  RECT 203.140 500.640 206.680 501.760 ;
  LAYER metal1 ;
  RECT 203.140 500.640 206.680 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 189.500 500.640 193.040 501.760 ;
  LAYER metal4 ;
  RECT 189.500 500.640 193.040 501.760 ;
  LAYER metal3 ;
  RECT 189.500 500.640 193.040 501.760 ;
  LAYER metal2 ;
  RECT 189.500 500.640 193.040 501.760 ;
  LAYER metal1 ;
  RECT 189.500 500.640 193.040 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 176.480 500.640 180.020 501.760 ;
  LAYER metal4 ;
  RECT 176.480 500.640 180.020 501.760 ;
  LAYER metal3 ;
  RECT 176.480 500.640 180.020 501.760 ;
  LAYER metal2 ;
  RECT 176.480 500.640 180.020 501.760 ;
  LAYER metal1 ;
  RECT 176.480 500.640 180.020 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 162.840 500.640 166.380 501.760 ;
  LAYER metal4 ;
  RECT 162.840 500.640 166.380 501.760 ;
  LAYER metal3 ;
  RECT 162.840 500.640 166.380 501.760 ;
  LAYER metal2 ;
  RECT 162.840 500.640 166.380 501.760 ;
  LAYER metal1 ;
  RECT 162.840 500.640 166.380 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 149.200 500.640 152.740 501.760 ;
  LAYER metal4 ;
  RECT 149.200 500.640 152.740 501.760 ;
  LAYER metal3 ;
  RECT 149.200 500.640 152.740 501.760 ;
  LAYER metal2 ;
  RECT 149.200 500.640 152.740 501.760 ;
  LAYER metal1 ;
  RECT 149.200 500.640 152.740 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 82.240 500.640 85.780 501.760 ;
  LAYER metal4 ;
  RECT 82.240 500.640 85.780 501.760 ;
  LAYER metal3 ;
  RECT 82.240 500.640 85.780 501.760 ;
  LAYER metal2 ;
  RECT 82.240 500.640 85.780 501.760 ;
  LAYER metal1 ;
  RECT 82.240 500.640 85.780 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 68.600 500.640 72.140 501.760 ;
  LAYER metal4 ;
  RECT 68.600 500.640 72.140 501.760 ;
  LAYER metal3 ;
  RECT 68.600 500.640 72.140 501.760 ;
  LAYER metal2 ;
  RECT 68.600 500.640 72.140 501.760 ;
  LAYER metal1 ;
  RECT 68.600 500.640 72.140 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 54.960 500.640 58.500 501.760 ;
  LAYER metal4 ;
  RECT 54.960 500.640 58.500 501.760 ;
  LAYER metal3 ;
  RECT 54.960 500.640 58.500 501.760 ;
  LAYER metal2 ;
  RECT 54.960 500.640 58.500 501.760 ;
  LAYER metal1 ;
  RECT 54.960 500.640 58.500 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 41.940 500.640 45.480 501.760 ;
  LAYER metal4 ;
  RECT 41.940 500.640 45.480 501.760 ;
  LAYER metal3 ;
  RECT 41.940 500.640 45.480 501.760 ;
  LAYER metal2 ;
  RECT 41.940 500.640 45.480 501.760 ;
  LAYER metal1 ;
  RECT 41.940 500.640 45.480 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 28.300 500.640 31.840 501.760 ;
  LAYER metal4 ;
  RECT 28.300 500.640 31.840 501.760 ;
  LAYER metal3 ;
  RECT 28.300 500.640 31.840 501.760 ;
  LAYER metal2 ;
  RECT 28.300 500.640 31.840 501.760 ;
  LAYER metal1 ;
  RECT 28.300 500.640 31.840 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 14.660 500.640 18.200 501.760 ;
  LAYER metal4 ;
  RECT 14.660 500.640 18.200 501.760 ;
  LAYER metal3 ;
  RECT 14.660 500.640 18.200 501.760 ;
  LAYER metal2 ;
  RECT 14.660 500.640 18.200 501.760 ;
  LAYER metal1 ;
  RECT 14.660 500.640 18.200 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3579.660 0.000 3583.200 1.120 ;
  LAYER metal4 ;
  RECT 3579.660 0.000 3583.200 1.120 ;
  LAYER metal3 ;
  RECT 3579.660 0.000 3583.200 1.120 ;
  LAYER metal2 ;
  RECT 3579.660 0.000 3583.200 1.120 ;
  LAYER metal1 ;
  RECT 3579.660 0.000 3583.200 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3566.020 0.000 3569.560 1.120 ;
  LAYER metal4 ;
  RECT 3566.020 0.000 3569.560 1.120 ;
  LAYER metal3 ;
  RECT 3566.020 0.000 3569.560 1.120 ;
  LAYER metal2 ;
  RECT 3566.020 0.000 3569.560 1.120 ;
  LAYER metal1 ;
  RECT 3566.020 0.000 3569.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3553.000 0.000 3556.540 1.120 ;
  LAYER metal4 ;
  RECT 3553.000 0.000 3556.540 1.120 ;
  LAYER metal3 ;
  RECT 3553.000 0.000 3556.540 1.120 ;
  LAYER metal2 ;
  RECT 3553.000 0.000 3556.540 1.120 ;
  LAYER metal1 ;
  RECT 3553.000 0.000 3556.540 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3539.360 0.000 3542.900 1.120 ;
  LAYER metal4 ;
  RECT 3539.360 0.000 3542.900 1.120 ;
  LAYER metal3 ;
  RECT 3539.360 0.000 3542.900 1.120 ;
  LAYER metal2 ;
  RECT 3539.360 0.000 3542.900 1.120 ;
  LAYER metal1 ;
  RECT 3539.360 0.000 3542.900 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3525.720 0.000 3529.260 1.120 ;
  LAYER metal4 ;
  RECT 3525.720 0.000 3529.260 1.120 ;
  LAYER metal3 ;
  RECT 3525.720 0.000 3529.260 1.120 ;
  LAYER metal2 ;
  RECT 3525.720 0.000 3529.260 1.120 ;
  LAYER metal1 ;
  RECT 3525.720 0.000 3529.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3458.760 0.000 3462.300 1.120 ;
  LAYER metal4 ;
  RECT 3458.760 0.000 3462.300 1.120 ;
  LAYER metal3 ;
  RECT 3458.760 0.000 3462.300 1.120 ;
  LAYER metal2 ;
  RECT 3458.760 0.000 3462.300 1.120 ;
  LAYER metal1 ;
  RECT 3458.760 0.000 3462.300 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3445.120 0.000 3448.660 1.120 ;
  LAYER metal4 ;
  RECT 3445.120 0.000 3448.660 1.120 ;
  LAYER metal3 ;
  RECT 3445.120 0.000 3448.660 1.120 ;
  LAYER metal2 ;
  RECT 3445.120 0.000 3448.660 1.120 ;
  LAYER metal1 ;
  RECT 3445.120 0.000 3448.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3432.100 0.000 3435.640 1.120 ;
  LAYER metal4 ;
  RECT 3432.100 0.000 3435.640 1.120 ;
  LAYER metal3 ;
  RECT 3432.100 0.000 3435.640 1.120 ;
  LAYER metal2 ;
  RECT 3432.100 0.000 3435.640 1.120 ;
  LAYER metal1 ;
  RECT 3432.100 0.000 3435.640 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3418.460 0.000 3422.000 1.120 ;
  LAYER metal4 ;
  RECT 3418.460 0.000 3422.000 1.120 ;
  LAYER metal3 ;
  RECT 3418.460 0.000 3422.000 1.120 ;
  LAYER metal2 ;
  RECT 3418.460 0.000 3422.000 1.120 ;
  LAYER metal1 ;
  RECT 3418.460 0.000 3422.000 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3404.820 0.000 3408.360 1.120 ;
  LAYER metal4 ;
  RECT 3404.820 0.000 3408.360 1.120 ;
  LAYER metal3 ;
  RECT 3404.820 0.000 3408.360 1.120 ;
  LAYER metal2 ;
  RECT 3404.820 0.000 3408.360 1.120 ;
  LAYER metal1 ;
  RECT 3404.820 0.000 3408.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3391.800 0.000 3395.340 1.120 ;
  LAYER metal4 ;
  RECT 3391.800 0.000 3395.340 1.120 ;
  LAYER metal3 ;
  RECT 3391.800 0.000 3395.340 1.120 ;
  LAYER metal2 ;
  RECT 3391.800 0.000 3395.340 1.120 ;
  LAYER metal1 ;
  RECT 3391.800 0.000 3395.340 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3324.220 0.000 3327.760 1.120 ;
  LAYER metal4 ;
  RECT 3324.220 0.000 3327.760 1.120 ;
  LAYER metal3 ;
  RECT 3324.220 0.000 3327.760 1.120 ;
  LAYER metal2 ;
  RECT 3324.220 0.000 3327.760 1.120 ;
  LAYER metal1 ;
  RECT 3324.220 0.000 3327.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3311.200 0.000 3314.740 1.120 ;
  LAYER metal4 ;
  RECT 3311.200 0.000 3314.740 1.120 ;
  LAYER metal3 ;
  RECT 3311.200 0.000 3314.740 1.120 ;
  LAYER metal2 ;
  RECT 3311.200 0.000 3314.740 1.120 ;
  LAYER metal1 ;
  RECT 3311.200 0.000 3314.740 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3297.560 0.000 3301.100 1.120 ;
  LAYER metal4 ;
  RECT 3297.560 0.000 3301.100 1.120 ;
  LAYER metal3 ;
  RECT 3297.560 0.000 3301.100 1.120 ;
  LAYER metal2 ;
  RECT 3297.560 0.000 3301.100 1.120 ;
  LAYER metal1 ;
  RECT 3297.560 0.000 3301.100 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3283.920 0.000 3287.460 1.120 ;
  LAYER metal4 ;
  RECT 3283.920 0.000 3287.460 1.120 ;
  LAYER metal3 ;
  RECT 3283.920 0.000 3287.460 1.120 ;
  LAYER metal2 ;
  RECT 3283.920 0.000 3287.460 1.120 ;
  LAYER metal1 ;
  RECT 3283.920 0.000 3287.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3270.900 0.000 3274.440 1.120 ;
  LAYER metal4 ;
  RECT 3270.900 0.000 3274.440 1.120 ;
  LAYER metal3 ;
  RECT 3270.900 0.000 3274.440 1.120 ;
  LAYER metal2 ;
  RECT 3270.900 0.000 3274.440 1.120 ;
  LAYER metal1 ;
  RECT 3270.900 0.000 3274.440 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3257.260 0.000 3260.800 1.120 ;
  LAYER metal4 ;
  RECT 3257.260 0.000 3260.800 1.120 ;
  LAYER metal3 ;
  RECT 3257.260 0.000 3260.800 1.120 ;
  LAYER metal2 ;
  RECT 3257.260 0.000 3260.800 1.120 ;
  LAYER metal1 ;
  RECT 3257.260 0.000 3260.800 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3190.300 0.000 3193.840 1.120 ;
  LAYER metal4 ;
  RECT 3190.300 0.000 3193.840 1.120 ;
  LAYER metal3 ;
  RECT 3190.300 0.000 3193.840 1.120 ;
  LAYER metal2 ;
  RECT 3190.300 0.000 3193.840 1.120 ;
  LAYER metal1 ;
  RECT 3190.300 0.000 3193.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3176.660 0.000 3180.200 1.120 ;
  LAYER metal4 ;
  RECT 3176.660 0.000 3180.200 1.120 ;
  LAYER metal3 ;
  RECT 3176.660 0.000 3180.200 1.120 ;
  LAYER metal2 ;
  RECT 3176.660 0.000 3180.200 1.120 ;
  LAYER metal1 ;
  RECT 3176.660 0.000 3180.200 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3163.020 0.000 3166.560 1.120 ;
  LAYER metal4 ;
  RECT 3163.020 0.000 3166.560 1.120 ;
  LAYER metal3 ;
  RECT 3163.020 0.000 3166.560 1.120 ;
  LAYER metal2 ;
  RECT 3163.020 0.000 3166.560 1.120 ;
  LAYER metal1 ;
  RECT 3163.020 0.000 3166.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3149.380 0.000 3152.920 1.120 ;
  LAYER metal4 ;
  RECT 3149.380 0.000 3152.920 1.120 ;
  LAYER metal3 ;
  RECT 3149.380 0.000 3152.920 1.120 ;
  LAYER metal2 ;
  RECT 3149.380 0.000 3152.920 1.120 ;
  LAYER metal1 ;
  RECT 3149.380 0.000 3152.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3136.360 0.000 3139.900 1.120 ;
  LAYER metal4 ;
  RECT 3136.360 0.000 3139.900 1.120 ;
  LAYER metal3 ;
  RECT 3136.360 0.000 3139.900 1.120 ;
  LAYER metal2 ;
  RECT 3136.360 0.000 3139.900 1.120 ;
  LAYER metal1 ;
  RECT 3136.360 0.000 3139.900 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3122.720 0.000 3126.260 1.120 ;
  LAYER metal4 ;
  RECT 3122.720 0.000 3126.260 1.120 ;
  LAYER metal3 ;
  RECT 3122.720 0.000 3126.260 1.120 ;
  LAYER metal2 ;
  RECT 3122.720 0.000 3126.260 1.120 ;
  LAYER metal1 ;
  RECT 3122.720 0.000 3126.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3055.760 0.000 3059.300 1.120 ;
  LAYER metal4 ;
  RECT 3055.760 0.000 3059.300 1.120 ;
  LAYER metal3 ;
  RECT 3055.760 0.000 3059.300 1.120 ;
  LAYER metal2 ;
  RECT 3055.760 0.000 3059.300 1.120 ;
  LAYER metal1 ;
  RECT 3055.760 0.000 3059.300 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3042.120 0.000 3045.660 1.120 ;
  LAYER metal4 ;
  RECT 3042.120 0.000 3045.660 1.120 ;
  LAYER metal3 ;
  RECT 3042.120 0.000 3045.660 1.120 ;
  LAYER metal2 ;
  RECT 3042.120 0.000 3045.660 1.120 ;
  LAYER metal1 ;
  RECT 3042.120 0.000 3045.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3028.480 0.000 3032.020 1.120 ;
  LAYER metal4 ;
  RECT 3028.480 0.000 3032.020 1.120 ;
  LAYER metal3 ;
  RECT 3028.480 0.000 3032.020 1.120 ;
  LAYER metal2 ;
  RECT 3028.480 0.000 3032.020 1.120 ;
  LAYER metal1 ;
  RECT 3028.480 0.000 3032.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3015.460 0.000 3019.000 1.120 ;
  LAYER metal4 ;
  RECT 3015.460 0.000 3019.000 1.120 ;
  LAYER metal3 ;
  RECT 3015.460 0.000 3019.000 1.120 ;
  LAYER metal2 ;
  RECT 3015.460 0.000 3019.000 1.120 ;
  LAYER metal1 ;
  RECT 3015.460 0.000 3019.000 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3001.820 0.000 3005.360 1.120 ;
  LAYER metal4 ;
  RECT 3001.820 0.000 3005.360 1.120 ;
  LAYER metal3 ;
  RECT 3001.820 0.000 3005.360 1.120 ;
  LAYER metal2 ;
  RECT 3001.820 0.000 3005.360 1.120 ;
  LAYER metal1 ;
  RECT 3001.820 0.000 3005.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2988.180 0.000 2991.720 1.120 ;
  LAYER metal4 ;
  RECT 2988.180 0.000 2991.720 1.120 ;
  LAYER metal3 ;
  RECT 2988.180 0.000 2991.720 1.120 ;
  LAYER metal2 ;
  RECT 2988.180 0.000 2991.720 1.120 ;
  LAYER metal1 ;
  RECT 2988.180 0.000 2991.720 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2921.220 0.000 2924.760 1.120 ;
  LAYER metal4 ;
  RECT 2921.220 0.000 2924.760 1.120 ;
  LAYER metal3 ;
  RECT 2921.220 0.000 2924.760 1.120 ;
  LAYER metal2 ;
  RECT 2921.220 0.000 2924.760 1.120 ;
  LAYER metal1 ;
  RECT 2921.220 0.000 2924.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2907.580 0.000 2911.120 1.120 ;
  LAYER metal4 ;
  RECT 2907.580 0.000 2911.120 1.120 ;
  LAYER metal3 ;
  RECT 2907.580 0.000 2911.120 1.120 ;
  LAYER metal2 ;
  RECT 2907.580 0.000 2911.120 1.120 ;
  LAYER metal1 ;
  RECT 2907.580 0.000 2911.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2894.560 0.000 2898.100 1.120 ;
  LAYER metal4 ;
  RECT 2894.560 0.000 2898.100 1.120 ;
  LAYER metal3 ;
  RECT 2894.560 0.000 2898.100 1.120 ;
  LAYER metal2 ;
  RECT 2894.560 0.000 2898.100 1.120 ;
  LAYER metal1 ;
  RECT 2894.560 0.000 2898.100 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2880.920 0.000 2884.460 1.120 ;
  LAYER metal4 ;
  RECT 2880.920 0.000 2884.460 1.120 ;
  LAYER metal3 ;
  RECT 2880.920 0.000 2884.460 1.120 ;
  LAYER metal2 ;
  RECT 2880.920 0.000 2884.460 1.120 ;
  LAYER metal1 ;
  RECT 2880.920 0.000 2884.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2867.280 0.000 2870.820 1.120 ;
  LAYER metal4 ;
  RECT 2867.280 0.000 2870.820 1.120 ;
  LAYER metal3 ;
  RECT 2867.280 0.000 2870.820 1.120 ;
  LAYER metal2 ;
  RECT 2867.280 0.000 2870.820 1.120 ;
  LAYER metal1 ;
  RECT 2867.280 0.000 2870.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2854.260 0.000 2857.800 1.120 ;
  LAYER metal4 ;
  RECT 2854.260 0.000 2857.800 1.120 ;
  LAYER metal3 ;
  RECT 2854.260 0.000 2857.800 1.120 ;
  LAYER metal2 ;
  RECT 2854.260 0.000 2857.800 1.120 ;
  LAYER metal1 ;
  RECT 2854.260 0.000 2857.800 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2786.680 0.000 2790.220 1.120 ;
  LAYER metal4 ;
  RECT 2786.680 0.000 2790.220 1.120 ;
  LAYER metal3 ;
  RECT 2786.680 0.000 2790.220 1.120 ;
  LAYER metal2 ;
  RECT 2786.680 0.000 2790.220 1.120 ;
  LAYER metal1 ;
  RECT 2786.680 0.000 2790.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2773.660 0.000 2777.200 1.120 ;
  LAYER metal4 ;
  RECT 2773.660 0.000 2777.200 1.120 ;
  LAYER metal3 ;
  RECT 2773.660 0.000 2777.200 1.120 ;
  LAYER metal2 ;
  RECT 2773.660 0.000 2777.200 1.120 ;
  LAYER metal1 ;
  RECT 2773.660 0.000 2777.200 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2760.020 0.000 2763.560 1.120 ;
  LAYER metal4 ;
  RECT 2760.020 0.000 2763.560 1.120 ;
  LAYER metal3 ;
  RECT 2760.020 0.000 2763.560 1.120 ;
  LAYER metal2 ;
  RECT 2760.020 0.000 2763.560 1.120 ;
  LAYER metal1 ;
  RECT 2760.020 0.000 2763.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2746.380 0.000 2749.920 1.120 ;
  LAYER metal4 ;
  RECT 2746.380 0.000 2749.920 1.120 ;
  LAYER metal3 ;
  RECT 2746.380 0.000 2749.920 1.120 ;
  LAYER metal2 ;
  RECT 2746.380 0.000 2749.920 1.120 ;
  LAYER metal1 ;
  RECT 2746.380 0.000 2749.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2732.740 0.000 2736.280 1.120 ;
  LAYER metal4 ;
  RECT 2732.740 0.000 2736.280 1.120 ;
  LAYER metal3 ;
  RECT 2732.740 0.000 2736.280 1.120 ;
  LAYER metal2 ;
  RECT 2732.740 0.000 2736.280 1.120 ;
  LAYER metal1 ;
  RECT 2732.740 0.000 2736.280 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2719.720 0.000 2723.260 1.120 ;
  LAYER metal4 ;
  RECT 2719.720 0.000 2723.260 1.120 ;
  LAYER metal3 ;
  RECT 2719.720 0.000 2723.260 1.120 ;
  LAYER metal2 ;
  RECT 2719.720 0.000 2723.260 1.120 ;
  LAYER metal1 ;
  RECT 2719.720 0.000 2723.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2652.140 0.000 2655.680 1.120 ;
  LAYER metal4 ;
  RECT 2652.140 0.000 2655.680 1.120 ;
  LAYER metal3 ;
  RECT 2652.140 0.000 2655.680 1.120 ;
  LAYER metal2 ;
  RECT 2652.140 0.000 2655.680 1.120 ;
  LAYER metal1 ;
  RECT 2652.140 0.000 2655.680 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2639.120 0.000 2642.660 1.120 ;
  LAYER metal4 ;
  RECT 2639.120 0.000 2642.660 1.120 ;
  LAYER metal3 ;
  RECT 2639.120 0.000 2642.660 1.120 ;
  LAYER metal2 ;
  RECT 2639.120 0.000 2642.660 1.120 ;
  LAYER metal1 ;
  RECT 2639.120 0.000 2642.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2625.480 0.000 2629.020 1.120 ;
  LAYER metal4 ;
  RECT 2625.480 0.000 2629.020 1.120 ;
  LAYER metal3 ;
  RECT 2625.480 0.000 2629.020 1.120 ;
  LAYER metal2 ;
  RECT 2625.480 0.000 2629.020 1.120 ;
  LAYER metal1 ;
  RECT 2625.480 0.000 2629.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2611.840 0.000 2615.380 1.120 ;
  LAYER metal4 ;
  RECT 2611.840 0.000 2615.380 1.120 ;
  LAYER metal3 ;
  RECT 2611.840 0.000 2615.380 1.120 ;
  LAYER metal2 ;
  RECT 2611.840 0.000 2615.380 1.120 ;
  LAYER metal1 ;
  RECT 2611.840 0.000 2615.380 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2598.820 0.000 2602.360 1.120 ;
  LAYER metal4 ;
  RECT 2598.820 0.000 2602.360 1.120 ;
  LAYER metal3 ;
  RECT 2598.820 0.000 2602.360 1.120 ;
  LAYER metal2 ;
  RECT 2598.820 0.000 2602.360 1.120 ;
  LAYER metal1 ;
  RECT 2598.820 0.000 2602.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2585.180 0.000 2588.720 1.120 ;
  LAYER metal4 ;
  RECT 2585.180 0.000 2588.720 1.120 ;
  LAYER metal3 ;
  RECT 2585.180 0.000 2588.720 1.120 ;
  LAYER metal2 ;
  RECT 2585.180 0.000 2588.720 1.120 ;
  LAYER metal1 ;
  RECT 2585.180 0.000 2588.720 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2518.220 0.000 2521.760 1.120 ;
  LAYER metal4 ;
  RECT 2518.220 0.000 2521.760 1.120 ;
  LAYER metal3 ;
  RECT 2518.220 0.000 2521.760 1.120 ;
  LAYER metal2 ;
  RECT 2518.220 0.000 2521.760 1.120 ;
  LAYER metal1 ;
  RECT 2518.220 0.000 2521.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2504.580 0.000 2508.120 1.120 ;
  LAYER metal4 ;
  RECT 2504.580 0.000 2508.120 1.120 ;
  LAYER metal3 ;
  RECT 2504.580 0.000 2508.120 1.120 ;
  LAYER metal2 ;
  RECT 2504.580 0.000 2508.120 1.120 ;
  LAYER metal1 ;
  RECT 2504.580 0.000 2508.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2490.940 0.000 2494.480 1.120 ;
  LAYER metal4 ;
  RECT 2490.940 0.000 2494.480 1.120 ;
  LAYER metal3 ;
  RECT 2490.940 0.000 2494.480 1.120 ;
  LAYER metal2 ;
  RECT 2490.940 0.000 2494.480 1.120 ;
  LAYER metal1 ;
  RECT 2490.940 0.000 2494.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2477.920 0.000 2481.460 1.120 ;
  LAYER metal4 ;
  RECT 2477.920 0.000 2481.460 1.120 ;
  LAYER metal3 ;
  RECT 2477.920 0.000 2481.460 1.120 ;
  LAYER metal2 ;
  RECT 2477.920 0.000 2481.460 1.120 ;
  LAYER metal1 ;
  RECT 2477.920 0.000 2481.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2464.280 0.000 2467.820 1.120 ;
  LAYER metal4 ;
  RECT 2464.280 0.000 2467.820 1.120 ;
  LAYER metal3 ;
  RECT 2464.280 0.000 2467.820 1.120 ;
  LAYER metal2 ;
  RECT 2464.280 0.000 2467.820 1.120 ;
  LAYER metal1 ;
  RECT 2464.280 0.000 2467.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2450.640 0.000 2454.180 1.120 ;
  LAYER metal4 ;
  RECT 2450.640 0.000 2454.180 1.120 ;
  LAYER metal3 ;
  RECT 2450.640 0.000 2454.180 1.120 ;
  LAYER metal2 ;
  RECT 2450.640 0.000 2454.180 1.120 ;
  LAYER metal1 ;
  RECT 2450.640 0.000 2454.180 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2383.680 0.000 2387.220 1.120 ;
  LAYER metal4 ;
  RECT 2383.680 0.000 2387.220 1.120 ;
  LAYER metal3 ;
  RECT 2383.680 0.000 2387.220 1.120 ;
  LAYER metal2 ;
  RECT 2383.680 0.000 2387.220 1.120 ;
  LAYER metal1 ;
  RECT 2383.680 0.000 2387.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2370.040 0.000 2373.580 1.120 ;
  LAYER metal4 ;
  RECT 2370.040 0.000 2373.580 1.120 ;
  LAYER metal3 ;
  RECT 2370.040 0.000 2373.580 1.120 ;
  LAYER metal2 ;
  RECT 2370.040 0.000 2373.580 1.120 ;
  LAYER metal1 ;
  RECT 2370.040 0.000 2373.580 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2357.020 0.000 2360.560 1.120 ;
  LAYER metal4 ;
  RECT 2357.020 0.000 2360.560 1.120 ;
  LAYER metal3 ;
  RECT 2357.020 0.000 2360.560 1.120 ;
  LAYER metal2 ;
  RECT 2357.020 0.000 2360.560 1.120 ;
  LAYER metal1 ;
  RECT 2357.020 0.000 2360.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2343.380 0.000 2346.920 1.120 ;
  LAYER metal4 ;
  RECT 2343.380 0.000 2346.920 1.120 ;
  LAYER metal3 ;
  RECT 2343.380 0.000 2346.920 1.120 ;
  LAYER metal2 ;
  RECT 2343.380 0.000 2346.920 1.120 ;
  LAYER metal1 ;
  RECT 2343.380 0.000 2346.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2329.740 0.000 2333.280 1.120 ;
  LAYER metal4 ;
  RECT 2329.740 0.000 2333.280 1.120 ;
  LAYER metal3 ;
  RECT 2329.740 0.000 2333.280 1.120 ;
  LAYER metal2 ;
  RECT 2329.740 0.000 2333.280 1.120 ;
  LAYER metal1 ;
  RECT 2329.740 0.000 2333.280 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2316.100 0.000 2319.640 1.120 ;
  LAYER metal4 ;
  RECT 2316.100 0.000 2319.640 1.120 ;
  LAYER metal3 ;
  RECT 2316.100 0.000 2319.640 1.120 ;
  LAYER metal2 ;
  RECT 2316.100 0.000 2319.640 1.120 ;
  LAYER metal1 ;
  RECT 2316.100 0.000 2319.640 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2249.140 0.000 2252.680 1.120 ;
  LAYER metal4 ;
  RECT 2249.140 0.000 2252.680 1.120 ;
  LAYER metal3 ;
  RECT 2249.140 0.000 2252.680 1.120 ;
  LAYER metal2 ;
  RECT 2249.140 0.000 2252.680 1.120 ;
  LAYER metal1 ;
  RECT 2249.140 0.000 2252.680 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2235.500 0.000 2239.040 1.120 ;
  LAYER metal4 ;
  RECT 2235.500 0.000 2239.040 1.120 ;
  LAYER metal3 ;
  RECT 2235.500 0.000 2239.040 1.120 ;
  LAYER metal2 ;
  RECT 2235.500 0.000 2239.040 1.120 ;
  LAYER metal1 ;
  RECT 2235.500 0.000 2239.040 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2222.480 0.000 2226.020 1.120 ;
  LAYER metal4 ;
  RECT 2222.480 0.000 2226.020 1.120 ;
  LAYER metal3 ;
  RECT 2222.480 0.000 2226.020 1.120 ;
  LAYER metal2 ;
  RECT 2222.480 0.000 2226.020 1.120 ;
  LAYER metal1 ;
  RECT 2222.480 0.000 2226.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2208.840 0.000 2212.380 1.120 ;
  LAYER metal4 ;
  RECT 2208.840 0.000 2212.380 1.120 ;
  LAYER metal3 ;
  RECT 2208.840 0.000 2212.380 1.120 ;
  LAYER metal2 ;
  RECT 2208.840 0.000 2212.380 1.120 ;
  LAYER metal1 ;
  RECT 2208.840 0.000 2212.380 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2195.200 0.000 2198.740 1.120 ;
  LAYER metal4 ;
  RECT 2195.200 0.000 2198.740 1.120 ;
  LAYER metal3 ;
  RECT 2195.200 0.000 2198.740 1.120 ;
  LAYER metal2 ;
  RECT 2195.200 0.000 2198.740 1.120 ;
  LAYER metal1 ;
  RECT 2195.200 0.000 2198.740 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2182.180 0.000 2185.720 1.120 ;
  LAYER metal4 ;
  RECT 2182.180 0.000 2185.720 1.120 ;
  LAYER metal3 ;
  RECT 2182.180 0.000 2185.720 1.120 ;
  LAYER metal2 ;
  RECT 2182.180 0.000 2185.720 1.120 ;
  LAYER metal1 ;
  RECT 2182.180 0.000 2185.720 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2114.600 0.000 2118.140 1.120 ;
  LAYER metal4 ;
  RECT 2114.600 0.000 2118.140 1.120 ;
  LAYER metal3 ;
  RECT 2114.600 0.000 2118.140 1.120 ;
  LAYER metal2 ;
  RECT 2114.600 0.000 2118.140 1.120 ;
  LAYER metal1 ;
  RECT 2114.600 0.000 2118.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2101.580 0.000 2105.120 1.120 ;
  LAYER metal4 ;
  RECT 2101.580 0.000 2105.120 1.120 ;
  LAYER metal3 ;
  RECT 2101.580 0.000 2105.120 1.120 ;
  LAYER metal2 ;
  RECT 2101.580 0.000 2105.120 1.120 ;
  LAYER metal1 ;
  RECT 2101.580 0.000 2105.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2087.940 0.000 2091.480 1.120 ;
  LAYER metal4 ;
  RECT 2087.940 0.000 2091.480 1.120 ;
  LAYER metal3 ;
  RECT 2087.940 0.000 2091.480 1.120 ;
  LAYER metal2 ;
  RECT 2087.940 0.000 2091.480 1.120 ;
  LAYER metal1 ;
  RECT 2087.940 0.000 2091.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2074.300 0.000 2077.840 1.120 ;
  LAYER metal4 ;
  RECT 2074.300 0.000 2077.840 1.120 ;
  LAYER metal3 ;
  RECT 2074.300 0.000 2077.840 1.120 ;
  LAYER metal2 ;
  RECT 2074.300 0.000 2077.840 1.120 ;
  LAYER metal1 ;
  RECT 2074.300 0.000 2077.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2061.280 0.000 2064.820 1.120 ;
  LAYER metal4 ;
  RECT 2061.280 0.000 2064.820 1.120 ;
  LAYER metal3 ;
  RECT 2061.280 0.000 2064.820 1.120 ;
  LAYER metal2 ;
  RECT 2061.280 0.000 2064.820 1.120 ;
  LAYER metal1 ;
  RECT 2061.280 0.000 2064.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2047.640 0.000 2051.180 1.120 ;
  LAYER metal4 ;
  RECT 2047.640 0.000 2051.180 1.120 ;
  LAYER metal3 ;
  RECT 2047.640 0.000 2051.180 1.120 ;
  LAYER metal2 ;
  RECT 2047.640 0.000 2051.180 1.120 ;
  LAYER metal1 ;
  RECT 2047.640 0.000 2051.180 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1980.680 0.000 1984.220 1.120 ;
  LAYER metal4 ;
  RECT 1980.680 0.000 1984.220 1.120 ;
  LAYER metal3 ;
  RECT 1980.680 0.000 1984.220 1.120 ;
  LAYER metal2 ;
  RECT 1980.680 0.000 1984.220 1.120 ;
  LAYER metal1 ;
  RECT 1980.680 0.000 1984.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1967.040 0.000 1970.580 1.120 ;
  LAYER metal4 ;
  RECT 1967.040 0.000 1970.580 1.120 ;
  LAYER metal3 ;
  RECT 1967.040 0.000 1970.580 1.120 ;
  LAYER metal2 ;
  RECT 1967.040 0.000 1970.580 1.120 ;
  LAYER metal1 ;
  RECT 1967.040 0.000 1970.580 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1953.400 0.000 1956.940 1.120 ;
  LAYER metal4 ;
  RECT 1953.400 0.000 1956.940 1.120 ;
  LAYER metal3 ;
  RECT 1953.400 0.000 1956.940 1.120 ;
  LAYER metal2 ;
  RECT 1953.400 0.000 1956.940 1.120 ;
  LAYER metal1 ;
  RECT 1953.400 0.000 1956.940 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1940.380 0.000 1943.920 1.120 ;
  LAYER metal4 ;
  RECT 1940.380 0.000 1943.920 1.120 ;
  LAYER metal3 ;
  RECT 1940.380 0.000 1943.920 1.120 ;
  LAYER metal2 ;
  RECT 1940.380 0.000 1943.920 1.120 ;
  LAYER metal1 ;
  RECT 1940.380 0.000 1943.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1926.740 0.000 1930.280 1.120 ;
  LAYER metal4 ;
  RECT 1926.740 0.000 1930.280 1.120 ;
  LAYER metal3 ;
  RECT 1926.740 0.000 1930.280 1.120 ;
  LAYER metal2 ;
  RECT 1926.740 0.000 1930.280 1.120 ;
  LAYER metal1 ;
  RECT 1926.740 0.000 1930.280 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1913.100 0.000 1916.640 1.120 ;
  LAYER metal4 ;
  RECT 1913.100 0.000 1916.640 1.120 ;
  LAYER metal3 ;
  RECT 1913.100 0.000 1916.640 1.120 ;
  LAYER metal2 ;
  RECT 1913.100 0.000 1916.640 1.120 ;
  LAYER metal1 ;
  RECT 1913.100 0.000 1916.640 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1850.480 0.000 1854.020 1.120 ;
  LAYER metal4 ;
  RECT 1850.480 0.000 1854.020 1.120 ;
  LAYER metal3 ;
  RECT 1850.480 0.000 1854.020 1.120 ;
  LAYER metal2 ;
  RECT 1850.480 0.000 1854.020 1.120 ;
  LAYER metal1 ;
  RECT 1850.480 0.000 1854.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1841.800 0.000 1845.340 1.120 ;
  LAYER metal4 ;
  RECT 1841.800 0.000 1845.340 1.120 ;
  LAYER metal3 ;
  RECT 1841.800 0.000 1845.340 1.120 ;
  LAYER metal2 ;
  RECT 1841.800 0.000 1845.340 1.120 ;
  LAYER metal1 ;
  RECT 1841.800 0.000 1845.340 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1828.780 0.000 1832.320 1.120 ;
  LAYER metal4 ;
  RECT 1828.780 0.000 1832.320 1.120 ;
  LAYER metal3 ;
  RECT 1828.780 0.000 1832.320 1.120 ;
  LAYER metal2 ;
  RECT 1828.780 0.000 1832.320 1.120 ;
  LAYER metal1 ;
  RECT 1828.780 0.000 1832.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1784.140 0.000 1787.680 1.120 ;
  LAYER metal4 ;
  RECT 1784.140 0.000 1787.680 1.120 ;
  LAYER metal3 ;
  RECT 1784.140 0.000 1787.680 1.120 ;
  LAYER metal2 ;
  RECT 1784.140 0.000 1787.680 1.120 ;
  LAYER metal1 ;
  RECT 1784.140 0.000 1787.680 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1761.200 0.000 1764.740 1.120 ;
  LAYER metal4 ;
  RECT 1761.200 0.000 1764.740 1.120 ;
  LAYER metal3 ;
  RECT 1761.200 0.000 1764.740 1.120 ;
  LAYER metal2 ;
  RECT 1761.200 0.000 1764.740 1.120 ;
  LAYER metal1 ;
  RECT 1761.200 0.000 1764.740 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1752.520 0.000 1756.060 1.120 ;
  LAYER metal4 ;
  RECT 1752.520 0.000 1756.060 1.120 ;
  LAYER metal3 ;
  RECT 1752.520 0.000 1756.060 1.120 ;
  LAYER metal2 ;
  RECT 1752.520 0.000 1756.060 1.120 ;
  LAYER metal1 ;
  RECT 1752.520 0.000 1756.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1694.860 0.000 1698.400 1.120 ;
  LAYER metal4 ;
  RECT 1694.860 0.000 1698.400 1.120 ;
  LAYER metal3 ;
  RECT 1694.860 0.000 1698.400 1.120 ;
  LAYER metal2 ;
  RECT 1694.860 0.000 1698.400 1.120 ;
  LAYER metal1 ;
  RECT 1694.860 0.000 1698.400 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1681.220 0.000 1684.760 1.120 ;
  LAYER metal4 ;
  RECT 1681.220 0.000 1684.760 1.120 ;
  LAYER metal3 ;
  RECT 1681.220 0.000 1684.760 1.120 ;
  LAYER metal2 ;
  RECT 1681.220 0.000 1684.760 1.120 ;
  LAYER metal1 ;
  RECT 1681.220 0.000 1684.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1668.200 0.000 1671.740 1.120 ;
  LAYER metal4 ;
  RECT 1668.200 0.000 1671.740 1.120 ;
  LAYER metal3 ;
  RECT 1668.200 0.000 1671.740 1.120 ;
  LAYER metal2 ;
  RECT 1668.200 0.000 1671.740 1.120 ;
  LAYER metal1 ;
  RECT 1668.200 0.000 1671.740 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1654.560 0.000 1658.100 1.120 ;
  LAYER metal4 ;
  RECT 1654.560 0.000 1658.100 1.120 ;
  LAYER metal3 ;
  RECT 1654.560 0.000 1658.100 1.120 ;
  LAYER metal2 ;
  RECT 1654.560 0.000 1658.100 1.120 ;
  LAYER metal1 ;
  RECT 1654.560 0.000 1658.100 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1640.920 0.000 1644.460 1.120 ;
  LAYER metal4 ;
  RECT 1640.920 0.000 1644.460 1.120 ;
  LAYER metal3 ;
  RECT 1640.920 0.000 1644.460 1.120 ;
  LAYER metal2 ;
  RECT 1640.920 0.000 1644.460 1.120 ;
  LAYER metal1 ;
  RECT 1640.920 0.000 1644.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1627.900 0.000 1631.440 1.120 ;
  LAYER metal4 ;
  RECT 1627.900 0.000 1631.440 1.120 ;
  LAYER metal3 ;
  RECT 1627.900 0.000 1631.440 1.120 ;
  LAYER metal2 ;
  RECT 1627.900 0.000 1631.440 1.120 ;
  LAYER metal1 ;
  RECT 1627.900 0.000 1631.440 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1560.320 0.000 1563.860 1.120 ;
  LAYER metal4 ;
  RECT 1560.320 0.000 1563.860 1.120 ;
  LAYER metal3 ;
  RECT 1560.320 0.000 1563.860 1.120 ;
  LAYER metal2 ;
  RECT 1560.320 0.000 1563.860 1.120 ;
  LAYER metal1 ;
  RECT 1560.320 0.000 1563.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1547.300 0.000 1550.840 1.120 ;
  LAYER metal4 ;
  RECT 1547.300 0.000 1550.840 1.120 ;
  LAYER metal3 ;
  RECT 1547.300 0.000 1550.840 1.120 ;
  LAYER metal2 ;
  RECT 1547.300 0.000 1550.840 1.120 ;
  LAYER metal1 ;
  RECT 1547.300 0.000 1550.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1533.660 0.000 1537.200 1.120 ;
  LAYER metal4 ;
  RECT 1533.660 0.000 1537.200 1.120 ;
  LAYER metal3 ;
  RECT 1533.660 0.000 1537.200 1.120 ;
  LAYER metal2 ;
  RECT 1533.660 0.000 1537.200 1.120 ;
  LAYER metal1 ;
  RECT 1533.660 0.000 1537.200 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1520.020 0.000 1523.560 1.120 ;
  LAYER metal4 ;
  RECT 1520.020 0.000 1523.560 1.120 ;
  LAYER metal3 ;
  RECT 1520.020 0.000 1523.560 1.120 ;
  LAYER metal2 ;
  RECT 1520.020 0.000 1523.560 1.120 ;
  LAYER metal1 ;
  RECT 1520.020 0.000 1523.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1507.000 0.000 1510.540 1.120 ;
  LAYER metal4 ;
  RECT 1507.000 0.000 1510.540 1.120 ;
  LAYER metal3 ;
  RECT 1507.000 0.000 1510.540 1.120 ;
  LAYER metal2 ;
  RECT 1507.000 0.000 1510.540 1.120 ;
  LAYER metal1 ;
  RECT 1507.000 0.000 1510.540 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1493.360 0.000 1496.900 1.120 ;
  LAYER metal4 ;
  RECT 1493.360 0.000 1496.900 1.120 ;
  LAYER metal3 ;
  RECT 1493.360 0.000 1496.900 1.120 ;
  LAYER metal2 ;
  RECT 1493.360 0.000 1496.900 1.120 ;
  LAYER metal1 ;
  RECT 1493.360 0.000 1496.900 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1426.400 0.000 1429.940 1.120 ;
  LAYER metal4 ;
  RECT 1426.400 0.000 1429.940 1.120 ;
  LAYER metal3 ;
  RECT 1426.400 0.000 1429.940 1.120 ;
  LAYER metal2 ;
  RECT 1426.400 0.000 1429.940 1.120 ;
  LAYER metal1 ;
  RECT 1426.400 0.000 1429.940 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1412.760 0.000 1416.300 1.120 ;
  LAYER metal4 ;
  RECT 1412.760 0.000 1416.300 1.120 ;
  LAYER metal3 ;
  RECT 1412.760 0.000 1416.300 1.120 ;
  LAYER metal2 ;
  RECT 1412.760 0.000 1416.300 1.120 ;
  LAYER metal1 ;
  RECT 1412.760 0.000 1416.300 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1399.120 0.000 1402.660 1.120 ;
  LAYER metal4 ;
  RECT 1399.120 0.000 1402.660 1.120 ;
  LAYER metal3 ;
  RECT 1399.120 0.000 1402.660 1.120 ;
  LAYER metal2 ;
  RECT 1399.120 0.000 1402.660 1.120 ;
  LAYER metal1 ;
  RECT 1399.120 0.000 1402.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1386.100 0.000 1389.640 1.120 ;
  LAYER metal4 ;
  RECT 1386.100 0.000 1389.640 1.120 ;
  LAYER metal3 ;
  RECT 1386.100 0.000 1389.640 1.120 ;
  LAYER metal2 ;
  RECT 1386.100 0.000 1389.640 1.120 ;
  LAYER metal1 ;
  RECT 1386.100 0.000 1389.640 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1372.460 0.000 1376.000 1.120 ;
  LAYER metal4 ;
  RECT 1372.460 0.000 1376.000 1.120 ;
  LAYER metal3 ;
  RECT 1372.460 0.000 1376.000 1.120 ;
  LAYER metal2 ;
  RECT 1372.460 0.000 1376.000 1.120 ;
  LAYER metal1 ;
  RECT 1372.460 0.000 1376.000 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1358.820 0.000 1362.360 1.120 ;
  LAYER metal4 ;
  RECT 1358.820 0.000 1362.360 1.120 ;
  LAYER metal3 ;
  RECT 1358.820 0.000 1362.360 1.120 ;
  LAYER metal2 ;
  RECT 1358.820 0.000 1362.360 1.120 ;
  LAYER metal1 ;
  RECT 1358.820 0.000 1362.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1291.860 0.000 1295.400 1.120 ;
  LAYER metal4 ;
  RECT 1291.860 0.000 1295.400 1.120 ;
  LAYER metal3 ;
  RECT 1291.860 0.000 1295.400 1.120 ;
  LAYER metal2 ;
  RECT 1291.860 0.000 1295.400 1.120 ;
  LAYER metal1 ;
  RECT 1291.860 0.000 1295.400 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1278.220 0.000 1281.760 1.120 ;
  LAYER metal4 ;
  RECT 1278.220 0.000 1281.760 1.120 ;
  LAYER metal3 ;
  RECT 1278.220 0.000 1281.760 1.120 ;
  LAYER metal2 ;
  RECT 1278.220 0.000 1281.760 1.120 ;
  LAYER metal1 ;
  RECT 1278.220 0.000 1281.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1264.580 0.000 1268.120 1.120 ;
  LAYER metal4 ;
  RECT 1264.580 0.000 1268.120 1.120 ;
  LAYER metal3 ;
  RECT 1264.580 0.000 1268.120 1.120 ;
  LAYER metal2 ;
  RECT 1264.580 0.000 1268.120 1.120 ;
  LAYER metal1 ;
  RECT 1264.580 0.000 1268.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1251.560 0.000 1255.100 1.120 ;
  LAYER metal4 ;
  RECT 1251.560 0.000 1255.100 1.120 ;
  LAYER metal3 ;
  RECT 1251.560 0.000 1255.100 1.120 ;
  LAYER metal2 ;
  RECT 1251.560 0.000 1255.100 1.120 ;
  LAYER metal1 ;
  RECT 1251.560 0.000 1255.100 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1237.920 0.000 1241.460 1.120 ;
  LAYER metal4 ;
  RECT 1237.920 0.000 1241.460 1.120 ;
  LAYER metal3 ;
  RECT 1237.920 0.000 1241.460 1.120 ;
  LAYER metal2 ;
  RECT 1237.920 0.000 1241.460 1.120 ;
  LAYER metal1 ;
  RECT 1237.920 0.000 1241.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1224.280 0.000 1227.820 1.120 ;
  LAYER metal4 ;
  RECT 1224.280 0.000 1227.820 1.120 ;
  LAYER metal3 ;
  RECT 1224.280 0.000 1227.820 1.120 ;
  LAYER metal2 ;
  RECT 1224.280 0.000 1227.820 1.120 ;
  LAYER metal1 ;
  RECT 1224.280 0.000 1227.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1157.320 0.000 1160.860 1.120 ;
  LAYER metal4 ;
  RECT 1157.320 0.000 1160.860 1.120 ;
  LAYER metal3 ;
  RECT 1157.320 0.000 1160.860 1.120 ;
  LAYER metal2 ;
  RECT 1157.320 0.000 1160.860 1.120 ;
  LAYER metal1 ;
  RECT 1157.320 0.000 1160.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1143.680 0.000 1147.220 1.120 ;
  LAYER metal4 ;
  RECT 1143.680 0.000 1147.220 1.120 ;
  LAYER metal3 ;
  RECT 1143.680 0.000 1147.220 1.120 ;
  LAYER metal2 ;
  RECT 1143.680 0.000 1147.220 1.120 ;
  LAYER metal1 ;
  RECT 1143.680 0.000 1147.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1130.660 0.000 1134.200 1.120 ;
  LAYER metal4 ;
  RECT 1130.660 0.000 1134.200 1.120 ;
  LAYER metal3 ;
  RECT 1130.660 0.000 1134.200 1.120 ;
  LAYER metal2 ;
  RECT 1130.660 0.000 1134.200 1.120 ;
  LAYER metal1 ;
  RECT 1130.660 0.000 1134.200 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1117.020 0.000 1120.560 1.120 ;
  LAYER metal4 ;
  RECT 1117.020 0.000 1120.560 1.120 ;
  LAYER metal3 ;
  RECT 1117.020 0.000 1120.560 1.120 ;
  LAYER metal2 ;
  RECT 1117.020 0.000 1120.560 1.120 ;
  LAYER metal1 ;
  RECT 1117.020 0.000 1120.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1103.380 0.000 1106.920 1.120 ;
  LAYER metal4 ;
  RECT 1103.380 0.000 1106.920 1.120 ;
  LAYER metal3 ;
  RECT 1103.380 0.000 1106.920 1.120 ;
  LAYER metal2 ;
  RECT 1103.380 0.000 1106.920 1.120 ;
  LAYER metal1 ;
  RECT 1103.380 0.000 1106.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1090.360 0.000 1093.900 1.120 ;
  LAYER metal4 ;
  RECT 1090.360 0.000 1093.900 1.120 ;
  LAYER metal3 ;
  RECT 1090.360 0.000 1093.900 1.120 ;
  LAYER metal2 ;
  RECT 1090.360 0.000 1093.900 1.120 ;
  LAYER metal1 ;
  RECT 1090.360 0.000 1093.900 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1022.780 0.000 1026.320 1.120 ;
  LAYER metal4 ;
  RECT 1022.780 0.000 1026.320 1.120 ;
  LAYER metal3 ;
  RECT 1022.780 0.000 1026.320 1.120 ;
  LAYER metal2 ;
  RECT 1022.780 0.000 1026.320 1.120 ;
  LAYER metal1 ;
  RECT 1022.780 0.000 1026.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1009.760 0.000 1013.300 1.120 ;
  LAYER metal4 ;
  RECT 1009.760 0.000 1013.300 1.120 ;
  LAYER metal3 ;
  RECT 1009.760 0.000 1013.300 1.120 ;
  LAYER metal2 ;
  RECT 1009.760 0.000 1013.300 1.120 ;
  LAYER metal1 ;
  RECT 1009.760 0.000 1013.300 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 996.120 0.000 999.660 1.120 ;
  LAYER metal4 ;
  RECT 996.120 0.000 999.660 1.120 ;
  LAYER metal3 ;
  RECT 996.120 0.000 999.660 1.120 ;
  LAYER metal2 ;
  RECT 996.120 0.000 999.660 1.120 ;
  LAYER metal1 ;
  RECT 996.120 0.000 999.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 982.480 0.000 986.020 1.120 ;
  LAYER metal4 ;
  RECT 982.480 0.000 986.020 1.120 ;
  LAYER metal3 ;
  RECT 982.480 0.000 986.020 1.120 ;
  LAYER metal2 ;
  RECT 982.480 0.000 986.020 1.120 ;
  LAYER metal1 ;
  RECT 982.480 0.000 986.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 969.460 0.000 973.000 1.120 ;
  LAYER metal4 ;
  RECT 969.460 0.000 973.000 1.120 ;
  LAYER metal3 ;
  RECT 969.460 0.000 973.000 1.120 ;
  LAYER metal2 ;
  RECT 969.460 0.000 973.000 1.120 ;
  LAYER metal1 ;
  RECT 969.460 0.000 973.000 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 955.820 0.000 959.360 1.120 ;
  LAYER metal4 ;
  RECT 955.820 0.000 959.360 1.120 ;
  LAYER metal3 ;
  RECT 955.820 0.000 959.360 1.120 ;
  LAYER metal2 ;
  RECT 955.820 0.000 959.360 1.120 ;
  LAYER metal1 ;
  RECT 955.820 0.000 959.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 888.240 0.000 891.780 1.120 ;
  LAYER metal4 ;
  RECT 888.240 0.000 891.780 1.120 ;
  LAYER metal3 ;
  RECT 888.240 0.000 891.780 1.120 ;
  LAYER metal2 ;
  RECT 888.240 0.000 891.780 1.120 ;
  LAYER metal1 ;
  RECT 888.240 0.000 891.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 875.220 0.000 878.760 1.120 ;
  LAYER metal4 ;
  RECT 875.220 0.000 878.760 1.120 ;
  LAYER metal3 ;
  RECT 875.220 0.000 878.760 1.120 ;
  LAYER metal2 ;
  RECT 875.220 0.000 878.760 1.120 ;
  LAYER metal1 ;
  RECT 875.220 0.000 878.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 861.580 0.000 865.120 1.120 ;
  LAYER metal4 ;
  RECT 861.580 0.000 865.120 1.120 ;
  LAYER metal3 ;
  RECT 861.580 0.000 865.120 1.120 ;
  LAYER metal2 ;
  RECT 861.580 0.000 865.120 1.120 ;
  LAYER metal1 ;
  RECT 861.580 0.000 865.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 847.940 0.000 851.480 1.120 ;
  LAYER metal4 ;
  RECT 847.940 0.000 851.480 1.120 ;
  LAYER metal3 ;
  RECT 847.940 0.000 851.480 1.120 ;
  LAYER metal2 ;
  RECT 847.940 0.000 851.480 1.120 ;
  LAYER metal1 ;
  RECT 847.940 0.000 851.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 834.920 0.000 838.460 1.120 ;
  LAYER metal4 ;
  RECT 834.920 0.000 838.460 1.120 ;
  LAYER metal3 ;
  RECT 834.920 0.000 838.460 1.120 ;
  LAYER metal2 ;
  RECT 834.920 0.000 838.460 1.120 ;
  LAYER metal1 ;
  RECT 834.920 0.000 838.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 821.280 0.000 824.820 1.120 ;
  LAYER metal4 ;
  RECT 821.280 0.000 824.820 1.120 ;
  LAYER metal3 ;
  RECT 821.280 0.000 824.820 1.120 ;
  LAYER metal2 ;
  RECT 821.280 0.000 824.820 1.120 ;
  LAYER metal1 ;
  RECT 821.280 0.000 824.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 754.320 0.000 757.860 1.120 ;
  LAYER metal4 ;
  RECT 754.320 0.000 757.860 1.120 ;
  LAYER metal3 ;
  RECT 754.320 0.000 757.860 1.120 ;
  LAYER metal2 ;
  RECT 754.320 0.000 757.860 1.120 ;
  LAYER metal1 ;
  RECT 754.320 0.000 757.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 740.680 0.000 744.220 1.120 ;
  LAYER metal4 ;
  RECT 740.680 0.000 744.220 1.120 ;
  LAYER metal3 ;
  RECT 740.680 0.000 744.220 1.120 ;
  LAYER metal2 ;
  RECT 740.680 0.000 744.220 1.120 ;
  LAYER metal1 ;
  RECT 740.680 0.000 744.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 727.040 0.000 730.580 1.120 ;
  LAYER metal4 ;
  RECT 727.040 0.000 730.580 1.120 ;
  LAYER metal3 ;
  RECT 727.040 0.000 730.580 1.120 ;
  LAYER metal2 ;
  RECT 727.040 0.000 730.580 1.120 ;
  LAYER metal1 ;
  RECT 727.040 0.000 730.580 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 714.020 0.000 717.560 1.120 ;
  LAYER metal4 ;
  RECT 714.020 0.000 717.560 1.120 ;
  LAYER metal3 ;
  RECT 714.020 0.000 717.560 1.120 ;
  LAYER metal2 ;
  RECT 714.020 0.000 717.560 1.120 ;
  LAYER metal1 ;
  RECT 714.020 0.000 717.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 700.380 0.000 703.920 1.120 ;
  LAYER metal4 ;
  RECT 700.380 0.000 703.920 1.120 ;
  LAYER metal3 ;
  RECT 700.380 0.000 703.920 1.120 ;
  LAYER metal2 ;
  RECT 700.380 0.000 703.920 1.120 ;
  LAYER metal1 ;
  RECT 700.380 0.000 703.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 686.740 0.000 690.280 1.120 ;
  LAYER metal4 ;
  RECT 686.740 0.000 690.280 1.120 ;
  LAYER metal3 ;
  RECT 686.740 0.000 690.280 1.120 ;
  LAYER metal2 ;
  RECT 686.740 0.000 690.280 1.120 ;
  LAYER metal1 ;
  RECT 686.740 0.000 690.280 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 619.780 0.000 623.320 1.120 ;
  LAYER metal4 ;
  RECT 619.780 0.000 623.320 1.120 ;
  LAYER metal3 ;
  RECT 619.780 0.000 623.320 1.120 ;
  LAYER metal2 ;
  RECT 619.780 0.000 623.320 1.120 ;
  LAYER metal1 ;
  RECT 619.780 0.000 623.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 606.140 0.000 609.680 1.120 ;
  LAYER metal4 ;
  RECT 606.140 0.000 609.680 1.120 ;
  LAYER metal3 ;
  RECT 606.140 0.000 609.680 1.120 ;
  LAYER metal2 ;
  RECT 606.140 0.000 609.680 1.120 ;
  LAYER metal1 ;
  RECT 606.140 0.000 609.680 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 593.120 0.000 596.660 1.120 ;
  LAYER metal4 ;
  RECT 593.120 0.000 596.660 1.120 ;
  LAYER metal3 ;
  RECT 593.120 0.000 596.660 1.120 ;
  LAYER metal2 ;
  RECT 593.120 0.000 596.660 1.120 ;
  LAYER metal1 ;
  RECT 593.120 0.000 596.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 579.480 0.000 583.020 1.120 ;
  LAYER metal4 ;
  RECT 579.480 0.000 583.020 1.120 ;
  LAYER metal3 ;
  RECT 579.480 0.000 583.020 1.120 ;
  LAYER metal2 ;
  RECT 579.480 0.000 583.020 1.120 ;
  LAYER metal1 ;
  RECT 579.480 0.000 583.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 565.840 0.000 569.380 1.120 ;
  LAYER metal4 ;
  RECT 565.840 0.000 569.380 1.120 ;
  LAYER metal3 ;
  RECT 565.840 0.000 569.380 1.120 ;
  LAYER metal2 ;
  RECT 565.840 0.000 569.380 1.120 ;
  LAYER metal1 ;
  RECT 565.840 0.000 569.380 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 552.820 0.000 556.360 1.120 ;
  LAYER metal4 ;
  RECT 552.820 0.000 556.360 1.120 ;
  LAYER metal3 ;
  RECT 552.820 0.000 556.360 1.120 ;
  LAYER metal2 ;
  RECT 552.820 0.000 556.360 1.120 ;
  LAYER metal1 ;
  RECT 552.820 0.000 556.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 485.240 0.000 488.780 1.120 ;
  LAYER metal4 ;
  RECT 485.240 0.000 488.780 1.120 ;
  LAYER metal3 ;
  RECT 485.240 0.000 488.780 1.120 ;
  LAYER metal2 ;
  RECT 485.240 0.000 488.780 1.120 ;
  LAYER metal1 ;
  RECT 485.240 0.000 488.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 471.600 0.000 475.140 1.120 ;
  LAYER metal4 ;
  RECT 471.600 0.000 475.140 1.120 ;
  LAYER metal3 ;
  RECT 471.600 0.000 475.140 1.120 ;
  LAYER metal2 ;
  RECT 471.600 0.000 475.140 1.120 ;
  LAYER metal1 ;
  RECT 471.600 0.000 475.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 458.580 0.000 462.120 1.120 ;
  LAYER metal4 ;
  RECT 458.580 0.000 462.120 1.120 ;
  LAYER metal3 ;
  RECT 458.580 0.000 462.120 1.120 ;
  LAYER metal2 ;
  RECT 458.580 0.000 462.120 1.120 ;
  LAYER metal1 ;
  RECT 458.580 0.000 462.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 444.940 0.000 448.480 1.120 ;
  LAYER metal4 ;
  RECT 444.940 0.000 448.480 1.120 ;
  LAYER metal3 ;
  RECT 444.940 0.000 448.480 1.120 ;
  LAYER metal2 ;
  RECT 444.940 0.000 448.480 1.120 ;
  LAYER metal1 ;
  RECT 444.940 0.000 448.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 431.300 0.000 434.840 1.120 ;
  LAYER metal4 ;
  RECT 431.300 0.000 434.840 1.120 ;
  LAYER metal3 ;
  RECT 431.300 0.000 434.840 1.120 ;
  LAYER metal2 ;
  RECT 431.300 0.000 434.840 1.120 ;
  LAYER metal1 ;
  RECT 431.300 0.000 434.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 418.280 0.000 421.820 1.120 ;
  LAYER metal4 ;
  RECT 418.280 0.000 421.820 1.120 ;
  LAYER metal3 ;
  RECT 418.280 0.000 421.820 1.120 ;
  LAYER metal2 ;
  RECT 418.280 0.000 421.820 1.120 ;
  LAYER metal1 ;
  RECT 418.280 0.000 421.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 350.700 0.000 354.240 1.120 ;
  LAYER metal4 ;
  RECT 350.700 0.000 354.240 1.120 ;
  LAYER metal3 ;
  RECT 350.700 0.000 354.240 1.120 ;
  LAYER metal2 ;
  RECT 350.700 0.000 354.240 1.120 ;
  LAYER metal1 ;
  RECT 350.700 0.000 354.240 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 337.680 0.000 341.220 1.120 ;
  LAYER metal4 ;
  RECT 337.680 0.000 341.220 1.120 ;
  LAYER metal3 ;
  RECT 337.680 0.000 341.220 1.120 ;
  LAYER metal2 ;
  RECT 337.680 0.000 341.220 1.120 ;
  LAYER metal1 ;
  RECT 337.680 0.000 341.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 324.040 0.000 327.580 1.120 ;
  LAYER metal4 ;
  RECT 324.040 0.000 327.580 1.120 ;
  LAYER metal3 ;
  RECT 324.040 0.000 327.580 1.120 ;
  LAYER metal2 ;
  RECT 324.040 0.000 327.580 1.120 ;
  LAYER metal1 ;
  RECT 324.040 0.000 327.580 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 310.400 0.000 313.940 1.120 ;
  LAYER metal4 ;
  RECT 310.400 0.000 313.940 1.120 ;
  LAYER metal3 ;
  RECT 310.400 0.000 313.940 1.120 ;
  LAYER metal2 ;
  RECT 310.400 0.000 313.940 1.120 ;
  LAYER metal1 ;
  RECT 310.400 0.000 313.940 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 297.380 0.000 300.920 1.120 ;
  LAYER metal4 ;
  RECT 297.380 0.000 300.920 1.120 ;
  LAYER metal3 ;
  RECT 297.380 0.000 300.920 1.120 ;
  LAYER metal2 ;
  RECT 297.380 0.000 300.920 1.120 ;
  LAYER metal1 ;
  RECT 297.380 0.000 300.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 283.740 0.000 287.280 1.120 ;
  LAYER metal4 ;
  RECT 283.740 0.000 287.280 1.120 ;
  LAYER metal3 ;
  RECT 283.740 0.000 287.280 1.120 ;
  LAYER metal2 ;
  RECT 283.740 0.000 287.280 1.120 ;
  LAYER metal1 ;
  RECT 283.740 0.000 287.280 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 216.780 0.000 220.320 1.120 ;
  LAYER metal4 ;
  RECT 216.780 0.000 220.320 1.120 ;
  LAYER metal3 ;
  RECT 216.780 0.000 220.320 1.120 ;
  LAYER metal2 ;
  RECT 216.780 0.000 220.320 1.120 ;
  LAYER metal1 ;
  RECT 216.780 0.000 220.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 203.140 0.000 206.680 1.120 ;
  LAYER metal4 ;
  RECT 203.140 0.000 206.680 1.120 ;
  LAYER metal3 ;
  RECT 203.140 0.000 206.680 1.120 ;
  LAYER metal2 ;
  RECT 203.140 0.000 206.680 1.120 ;
  LAYER metal1 ;
  RECT 203.140 0.000 206.680 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 189.500 0.000 193.040 1.120 ;
  LAYER metal4 ;
  RECT 189.500 0.000 193.040 1.120 ;
  LAYER metal3 ;
  RECT 189.500 0.000 193.040 1.120 ;
  LAYER metal2 ;
  RECT 189.500 0.000 193.040 1.120 ;
  LAYER metal1 ;
  RECT 189.500 0.000 193.040 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 176.480 0.000 180.020 1.120 ;
  LAYER metal4 ;
  RECT 176.480 0.000 180.020 1.120 ;
  LAYER metal3 ;
  RECT 176.480 0.000 180.020 1.120 ;
  LAYER metal2 ;
  RECT 176.480 0.000 180.020 1.120 ;
  LAYER metal1 ;
  RECT 176.480 0.000 180.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 162.840 0.000 166.380 1.120 ;
  LAYER metal4 ;
  RECT 162.840 0.000 166.380 1.120 ;
  LAYER metal3 ;
  RECT 162.840 0.000 166.380 1.120 ;
  LAYER metal2 ;
  RECT 162.840 0.000 166.380 1.120 ;
  LAYER metal1 ;
  RECT 162.840 0.000 166.380 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 149.200 0.000 152.740 1.120 ;
  LAYER metal4 ;
  RECT 149.200 0.000 152.740 1.120 ;
  LAYER metal3 ;
  RECT 149.200 0.000 152.740 1.120 ;
  LAYER metal2 ;
  RECT 149.200 0.000 152.740 1.120 ;
  LAYER metal1 ;
  RECT 149.200 0.000 152.740 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 82.240 0.000 85.780 1.120 ;
  LAYER metal4 ;
  RECT 82.240 0.000 85.780 1.120 ;
  LAYER metal3 ;
  RECT 82.240 0.000 85.780 1.120 ;
  LAYER metal2 ;
  RECT 82.240 0.000 85.780 1.120 ;
  LAYER metal1 ;
  RECT 82.240 0.000 85.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 68.600 0.000 72.140 1.120 ;
  LAYER metal4 ;
  RECT 68.600 0.000 72.140 1.120 ;
  LAYER metal3 ;
  RECT 68.600 0.000 72.140 1.120 ;
  LAYER metal2 ;
  RECT 68.600 0.000 72.140 1.120 ;
  LAYER metal1 ;
  RECT 68.600 0.000 72.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 54.960 0.000 58.500 1.120 ;
  LAYER metal4 ;
  RECT 54.960 0.000 58.500 1.120 ;
  LAYER metal3 ;
  RECT 54.960 0.000 58.500 1.120 ;
  LAYER metal2 ;
  RECT 54.960 0.000 58.500 1.120 ;
  LAYER metal1 ;
  RECT 54.960 0.000 58.500 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 41.940 0.000 45.480 1.120 ;
  LAYER metal4 ;
  RECT 41.940 0.000 45.480 1.120 ;
  LAYER metal3 ;
  RECT 41.940 0.000 45.480 1.120 ;
  LAYER metal2 ;
  RECT 41.940 0.000 45.480 1.120 ;
  LAYER metal1 ;
  RECT 41.940 0.000 45.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 28.300 0.000 31.840 1.120 ;
  LAYER metal4 ;
  RECT 28.300 0.000 31.840 1.120 ;
  LAYER metal3 ;
  RECT 28.300 0.000 31.840 1.120 ;
  LAYER metal2 ;
  RECT 28.300 0.000 31.840 1.120 ;
  LAYER metal1 ;
  RECT 28.300 0.000 31.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 14.660 0.000 18.200 1.120 ;
  LAYER metal4 ;
  RECT 14.660 0.000 18.200 1.120 ;
  LAYER metal3 ;
  RECT 14.660 0.000 18.200 1.120 ;
  LAYER metal2 ;
  RECT 14.660 0.000 18.200 1.120 ;
  LAYER metal1 ;
  RECT 14.660 0.000 18.200 1.120 ;
 END
END GND
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal5 ;
  RECT 3594.880 485.860 3596.000 489.100 ;
  LAYER metal4 ;
  RECT 3594.880 485.860 3596.000 489.100 ;
  LAYER metal3 ;
  RECT 3594.880 485.860 3596.000 489.100 ;
  LAYER metal2 ;
  RECT 3594.880 485.860 3596.000 489.100 ;
  LAYER metal1 ;
  RECT 3594.880 485.860 3596.000 489.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 478.020 3596.000 481.260 ;
  LAYER metal4 ;
  RECT 3594.880 478.020 3596.000 481.260 ;
  LAYER metal3 ;
  RECT 3594.880 478.020 3596.000 481.260 ;
  LAYER metal2 ;
  RECT 3594.880 478.020 3596.000 481.260 ;
  LAYER metal1 ;
  RECT 3594.880 478.020 3596.000 481.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 438.820 3596.000 442.060 ;
  LAYER metal4 ;
  RECT 3594.880 438.820 3596.000 442.060 ;
  LAYER metal3 ;
  RECT 3594.880 438.820 3596.000 442.060 ;
  LAYER metal2 ;
  RECT 3594.880 438.820 3596.000 442.060 ;
  LAYER metal1 ;
  RECT 3594.880 438.820 3596.000 442.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 430.980 3596.000 434.220 ;
  LAYER metal4 ;
  RECT 3594.880 430.980 3596.000 434.220 ;
  LAYER metal3 ;
  RECT 3594.880 430.980 3596.000 434.220 ;
  LAYER metal2 ;
  RECT 3594.880 430.980 3596.000 434.220 ;
  LAYER metal1 ;
  RECT 3594.880 430.980 3596.000 434.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 423.140 3596.000 426.380 ;
  LAYER metal4 ;
  RECT 3594.880 423.140 3596.000 426.380 ;
  LAYER metal3 ;
  RECT 3594.880 423.140 3596.000 426.380 ;
  LAYER metal2 ;
  RECT 3594.880 423.140 3596.000 426.380 ;
  LAYER metal1 ;
  RECT 3594.880 423.140 3596.000 426.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 415.300 3596.000 418.540 ;
  LAYER metal4 ;
  RECT 3594.880 415.300 3596.000 418.540 ;
  LAYER metal3 ;
  RECT 3594.880 415.300 3596.000 418.540 ;
  LAYER metal2 ;
  RECT 3594.880 415.300 3596.000 418.540 ;
  LAYER metal1 ;
  RECT 3594.880 415.300 3596.000 418.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 407.460 3596.000 410.700 ;
  LAYER metal4 ;
  RECT 3594.880 407.460 3596.000 410.700 ;
  LAYER metal3 ;
  RECT 3594.880 407.460 3596.000 410.700 ;
  LAYER metal2 ;
  RECT 3594.880 407.460 3596.000 410.700 ;
  LAYER metal1 ;
  RECT 3594.880 407.460 3596.000 410.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 399.620 3596.000 402.860 ;
  LAYER metal4 ;
  RECT 3594.880 399.620 3596.000 402.860 ;
  LAYER metal3 ;
  RECT 3594.880 399.620 3596.000 402.860 ;
  LAYER metal2 ;
  RECT 3594.880 399.620 3596.000 402.860 ;
  LAYER metal1 ;
  RECT 3594.880 399.620 3596.000 402.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 360.420 3596.000 363.660 ;
  LAYER metal4 ;
  RECT 3594.880 360.420 3596.000 363.660 ;
  LAYER metal3 ;
  RECT 3594.880 360.420 3596.000 363.660 ;
  LAYER metal2 ;
  RECT 3594.880 360.420 3596.000 363.660 ;
  LAYER metal1 ;
  RECT 3594.880 360.420 3596.000 363.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 352.580 3596.000 355.820 ;
  LAYER metal4 ;
  RECT 3594.880 352.580 3596.000 355.820 ;
  LAYER metal3 ;
  RECT 3594.880 352.580 3596.000 355.820 ;
  LAYER metal2 ;
  RECT 3594.880 352.580 3596.000 355.820 ;
  LAYER metal1 ;
  RECT 3594.880 352.580 3596.000 355.820 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 344.740 3596.000 347.980 ;
  LAYER metal4 ;
  RECT 3594.880 344.740 3596.000 347.980 ;
  LAYER metal3 ;
  RECT 3594.880 344.740 3596.000 347.980 ;
  LAYER metal2 ;
  RECT 3594.880 344.740 3596.000 347.980 ;
  LAYER metal1 ;
  RECT 3594.880 344.740 3596.000 347.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 336.900 3596.000 340.140 ;
  LAYER metal4 ;
  RECT 3594.880 336.900 3596.000 340.140 ;
  LAYER metal3 ;
  RECT 3594.880 336.900 3596.000 340.140 ;
  LAYER metal2 ;
  RECT 3594.880 336.900 3596.000 340.140 ;
  LAYER metal1 ;
  RECT 3594.880 336.900 3596.000 340.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 329.060 3596.000 332.300 ;
  LAYER metal4 ;
  RECT 3594.880 329.060 3596.000 332.300 ;
  LAYER metal3 ;
  RECT 3594.880 329.060 3596.000 332.300 ;
  LAYER metal2 ;
  RECT 3594.880 329.060 3596.000 332.300 ;
  LAYER metal1 ;
  RECT 3594.880 329.060 3596.000 332.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 321.220 3596.000 324.460 ;
  LAYER metal4 ;
  RECT 3594.880 321.220 3596.000 324.460 ;
  LAYER metal3 ;
  RECT 3594.880 321.220 3596.000 324.460 ;
  LAYER metal2 ;
  RECT 3594.880 321.220 3596.000 324.460 ;
  LAYER metal1 ;
  RECT 3594.880 321.220 3596.000 324.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 282.020 3596.000 285.260 ;
  LAYER metal4 ;
  RECT 3594.880 282.020 3596.000 285.260 ;
  LAYER metal3 ;
  RECT 3594.880 282.020 3596.000 285.260 ;
  LAYER metal2 ;
  RECT 3594.880 282.020 3596.000 285.260 ;
  LAYER metal1 ;
  RECT 3594.880 282.020 3596.000 285.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 274.180 3596.000 277.420 ;
  LAYER metal4 ;
  RECT 3594.880 274.180 3596.000 277.420 ;
  LAYER metal3 ;
  RECT 3594.880 274.180 3596.000 277.420 ;
  LAYER metal2 ;
  RECT 3594.880 274.180 3596.000 277.420 ;
  LAYER metal1 ;
  RECT 3594.880 274.180 3596.000 277.420 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 266.340 3596.000 269.580 ;
  LAYER metal4 ;
  RECT 3594.880 266.340 3596.000 269.580 ;
  LAYER metal3 ;
  RECT 3594.880 266.340 3596.000 269.580 ;
  LAYER metal2 ;
  RECT 3594.880 266.340 3596.000 269.580 ;
  LAYER metal1 ;
  RECT 3594.880 266.340 3596.000 269.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 258.500 3596.000 261.740 ;
  LAYER metal4 ;
  RECT 3594.880 258.500 3596.000 261.740 ;
  LAYER metal3 ;
  RECT 3594.880 258.500 3596.000 261.740 ;
  LAYER metal2 ;
  RECT 3594.880 258.500 3596.000 261.740 ;
  LAYER metal1 ;
  RECT 3594.880 258.500 3596.000 261.740 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 250.660 3596.000 253.900 ;
  LAYER metal4 ;
  RECT 3594.880 250.660 3596.000 253.900 ;
  LAYER metal3 ;
  RECT 3594.880 250.660 3596.000 253.900 ;
  LAYER metal2 ;
  RECT 3594.880 250.660 3596.000 253.900 ;
  LAYER metal1 ;
  RECT 3594.880 250.660 3596.000 253.900 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 242.820 3596.000 246.060 ;
  LAYER metal4 ;
  RECT 3594.880 242.820 3596.000 246.060 ;
  LAYER metal3 ;
  RECT 3594.880 242.820 3596.000 246.060 ;
  LAYER metal2 ;
  RECT 3594.880 242.820 3596.000 246.060 ;
  LAYER metal1 ;
  RECT 3594.880 242.820 3596.000 246.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 203.620 3596.000 206.860 ;
  LAYER metal4 ;
  RECT 3594.880 203.620 3596.000 206.860 ;
  LAYER metal3 ;
  RECT 3594.880 203.620 3596.000 206.860 ;
  LAYER metal2 ;
  RECT 3594.880 203.620 3596.000 206.860 ;
  LAYER metal1 ;
  RECT 3594.880 203.620 3596.000 206.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 195.780 3596.000 199.020 ;
  LAYER metal4 ;
  RECT 3594.880 195.780 3596.000 199.020 ;
  LAYER metal3 ;
  RECT 3594.880 195.780 3596.000 199.020 ;
  LAYER metal2 ;
  RECT 3594.880 195.780 3596.000 199.020 ;
  LAYER metal1 ;
  RECT 3594.880 195.780 3596.000 199.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 187.940 3596.000 191.180 ;
  LAYER metal4 ;
  RECT 3594.880 187.940 3596.000 191.180 ;
  LAYER metal3 ;
  RECT 3594.880 187.940 3596.000 191.180 ;
  LAYER metal2 ;
  RECT 3594.880 187.940 3596.000 191.180 ;
  LAYER metal1 ;
  RECT 3594.880 187.940 3596.000 191.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 180.100 3596.000 183.340 ;
  LAYER metal4 ;
  RECT 3594.880 180.100 3596.000 183.340 ;
  LAYER metal3 ;
  RECT 3594.880 180.100 3596.000 183.340 ;
  LAYER metal2 ;
  RECT 3594.880 180.100 3596.000 183.340 ;
  LAYER metal1 ;
  RECT 3594.880 180.100 3596.000 183.340 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 172.260 3596.000 175.500 ;
  LAYER metal4 ;
  RECT 3594.880 172.260 3596.000 175.500 ;
  LAYER metal3 ;
  RECT 3594.880 172.260 3596.000 175.500 ;
  LAYER metal2 ;
  RECT 3594.880 172.260 3596.000 175.500 ;
  LAYER metal1 ;
  RECT 3594.880 172.260 3596.000 175.500 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 164.420 3596.000 167.660 ;
  LAYER metal4 ;
  RECT 3594.880 164.420 3596.000 167.660 ;
  LAYER metal3 ;
  RECT 3594.880 164.420 3596.000 167.660 ;
  LAYER metal2 ;
  RECT 3594.880 164.420 3596.000 167.660 ;
  LAYER metal1 ;
  RECT 3594.880 164.420 3596.000 167.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 125.220 3596.000 128.460 ;
  LAYER metal4 ;
  RECT 3594.880 125.220 3596.000 128.460 ;
  LAYER metal3 ;
  RECT 3594.880 125.220 3596.000 128.460 ;
  LAYER metal2 ;
  RECT 3594.880 125.220 3596.000 128.460 ;
  LAYER metal1 ;
  RECT 3594.880 125.220 3596.000 128.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 117.380 3596.000 120.620 ;
  LAYER metal4 ;
  RECT 3594.880 117.380 3596.000 120.620 ;
  LAYER metal3 ;
  RECT 3594.880 117.380 3596.000 120.620 ;
  LAYER metal2 ;
  RECT 3594.880 117.380 3596.000 120.620 ;
  LAYER metal1 ;
  RECT 3594.880 117.380 3596.000 120.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 109.540 3596.000 112.780 ;
  LAYER metal4 ;
  RECT 3594.880 109.540 3596.000 112.780 ;
  LAYER metal3 ;
  RECT 3594.880 109.540 3596.000 112.780 ;
  LAYER metal2 ;
  RECT 3594.880 109.540 3596.000 112.780 ;
  LAYER metal1 ;
  RECT 3594.880 109.540 3596.000 112.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 101.700 3596.000 104.940 ;
  LAYER metal4 ;
  RECT 3594.880 101.700 3596.000 104.940 ;
  LAYER metal3 ;
  RECT 3594.880 101.700 3596.000 104.940 ;
  LAYER metal2 ;
  RECT 3594.880 101.700 3596.000 104.940 ;
  LAYER metal1 ;
  RECT 3594.880 101.700 3596.000 104.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 93.860 3596.000 97.100 ;
  LAYER metal4 ;
  RECT 3594.880 93.860 3596.000 97.100 ;
  LAYER metal3 ;
  RECT 3594.880 93.860 3596.000 97.100 ;
  LAYER metal2 ;
  RECT 3594.880 93.860 3596.000 97.100 ;
  LAYER metal1 ;
  RECT 3594.880 93.860 3596.000 97.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 86.020 3596.000 89.260 ;
  LAYER metal4 ;
  RECT 3594.880 86.020 3596.000 89.260 ;
  LAYER metal3 ;
  RECT 3594.880 86.020 3596.000 89.260 ;
  LAYER metal2 ;
  RECT 3594.880 86.020 3596.000 89.260 ;
  LAYER metal1 ;
  RECT 3594.880 86.020 3596.000 89.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 46.820 3596.000 50.060 ;
  LAYER metal4 ;
  RECT 3594.880 46.820 3596.000 50.060 ;
  LAYER metal3 ;
  RECT 3594.880 46.820 3596.000 50.060 ;
  LAYER metal2 ;
  RECT 3594.880 46.820 3596.000 50.060 ;
  LAYER metal1 ;
  RECT 3594.880 46.820 3596.000 50.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 38.980 3596.000 42.220 ;
  LAYER metal4 ;
  RECT 3594.880 38.980 3596.000 42.220 ;
  LAYER metal3 ;
  RECT 3594.880 38.980 3596.000 42.220 ;
  LAYER metal2 ;
  RECT 3594.880 38.980 3596.000 42.220 ;
  LAYER metal1 ;
  RECT 3594.880 38.980 3596.000 42.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 31.140 3596.000 34.380 ;
  LAYER metal4 ;
  RECT 3594.880 31.140 3596.000 34.380 ;
  LAYER metal3 ;
  RECT 3594.880 31.140 3596.000 34.380 ;
  LAYER metal2 ;
  RECT 3594.880 31.140 3596.000 34.380 ;
  LAYER metal1 ;
  RECT 3594.880 31.140 3596.000 34.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 23.300 3596.000 26.540 ;
  LAYER metal4 ;
  RECT 3594.880 23.300 3596.000 26.540 ;
  LAYER metal3 ;
  RECT 3594.880 23.300 3596.000 26.540 ;
  LAYER metal2 ;
  RECT 3594.880 23.300 3596.000 26.540 ;
  LAYER metal1 ;
  RECT 3594.880 23.300 3596.000 26.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 15.460 3596.000 18.700 ;
  LAYER metal4 ;
  RECT 3594.880 15.460 3596.000 18.700 ;
  LAYER metal3 ;
  RECT 3594.880 15.460 3596.000 18.700 ;
  LAYER metal2 ;
  RECT 3594.880 15.460 3596.000 18.700 ;
  LAYER metal1 ;
  RECT 3594.880 15.460 3596.000 18.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3594.880 7.620 3596.000 10.860 ;
  LAYER metal4 ;
  RECT 3594.880 7.620 3596.000 10.860 ;
  LAYER metal3 ;
  RECT 3594.880 7.620 3596.000 10.860 ;
  LAYER metal2 ;
  RECT 3594.880 7.620 3596.000 10.860 ;
  LAYER metal1 ;
  RECT 3594.880 7.620 3596.000 10.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 485.860 1.120 489.100 ;
  LAYER metal4 ;
  RECT 0.000 485.860 1.120 489.100 ;
  LAYER metal3 ;
  RECT 0.000 485.860 1.120 489.100 ;
  LAYER metal2 ;
  RECT 0.000 485.860 1.120 489.100 ;
  LAYER metal1 ;
  RECT 0.000 485.860 1.120 489.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 478.020 1.120 481.260 ;
  LAYER metal4 ;
  RECT 0.000 478.020 1.120 481.260 ;
  LAYER metal3 ;
  RECT 0.000 478.020 1.120 481.260 ;
  LAYER metal2 ;
  RECT 0.000 478.020 1.120 481.260 ;
  LAYER metal1 ;
  RECT 0.000 478.020 1.120 481.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 438.820 1.120 442.060 ;
  LAYER metal4 ;
  RECT 0.000 438.820 1.120 442.060 ;
  LAYER metal3 ;
  RECT 0.000 438.820 1.120 442.060 ;
  LAYER metal2 ;
  RECT 0.000 438.820 1.120 442.060 ;
  LAYER metal1 ;
  RECT 0.000 438.820 1.120 442.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 430.980 1.120 434.220 ;
  LAYER metal4 ;
  RECT 0.000 430.980 1.120 434.220 ;
  LAYER metal3 ;
  RECT 0.000 430.980 1.120 434.220 ;
  LAYER metal2 ;
  RECT 0.000 430.980 1.120 434.220 ;
  LAYER metal1 ;
  RECT 0.000 430.980 1.120 434.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 423.140 1.120 426.380 ;
  LAYER metal4 ;
  RECT 0.000 423.140 1.120 426.380 ;
  LAYER metal3 ;
  RECT 0.000 423.140 1.120 426.380 ;
  LAYER metal2 ;
  RECT 0.000 423.140 1.120 426.380 ;
  LAYER metal1 ;
  RECT 0.000 423.140 1.120 426.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 415.300 1.120 418.540 ;
  LAYER metal4 ;
  RECT 0.000 415.300 1.120 418.540 ;
  LAYER metal3 ;
  RECT 0.000 415.300 1.120 418.540 ;
  LAYER metal2 ;
  RECT 0.000 415.300 1.120 418.540 ;
  LAYER metal1 ;
  RECT 0.000 415.300 1.120 418.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 407.460 1.120 410.700 ;
  LAYER metal4 ;
  RECT 0.000 407.460 1.120 410.700 ;
  LAYER metal3 ;
  RECT 0.000 407.460 1.120 410.700 ;
  LAYER metal2 ;
  RECT 0.000 407.460 1.120 410.700 ;
  LAYER metal1 ;
  RECT 0.000 407.460 1.120 410.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 399.620 1.120 402.860 ;
  LAYER metal4 ;
  RECT 0.000 399.620 1.120 402.860 ;
  LAYER metal3 ;
  RECT 0.000 399.620 1.120 402.860 ;
  LAYER metal2 ;
  RECT 0.000 399.620 1.120 402.860 ;
  LAYER metal1 ;
  RECT 0.000 399.620 1.120 402.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 360.420 1.120 363.660 ;
  LAYER metal4 ;
  RECT 0.000 360.420 1.120 363.660 ;
  LAYER metal3 ;
  RECT 0.000 360.420 1.120 363.660 ;
  LAYER metal2 ;
  RECT 0.000 360.420 1.120 363.660 ;
  LAYER metal1 ;
  RECT 0.000 360.420 1.120 363.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 352.580 1.120 355.820 ;
  LAYER metal4 ;
  RECT 0.000 352.580 1.120 355.820 ;
  LAYER metal3 ;
  RECT 0.000 352.580 1.120 355.820 ;
  LAYER metal2 ;
  RECT 0.000 352.580 1.120 355.820 ;
  LAYER metal1 ;
  RECT 0.000 352.580 1.120 355.820 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 344.740 1.120 347.980 ;
  LAYER metal4 ;
  RECT 0.000 344.740 1.120 347.980 ;
  LAYER metal3 ;
  RECT 0.000 344.740 1.120 347.980 ;
  LAYER metal2 ;
  RECT 0.000 344.740 1.120 347.980 ;
  LAYER metal1 ;
  RECT 0.000 344.740 1.120 347.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 336.900 1.120 340.140 ;
  LAYER metal4 ;
  RECT 0.000 336.900 1.120 340.140 ;
  LAYER metal3 ;
  RECT 0.000 336.900 1.120 340.140 ;
  LAYER metal2 ;
  RECT 0.000 336.900 1.120 340.140 ;
  LAYER metal1 ;
  RECT 0.000 336.900 1.120 340.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 329.060 1.120 332.300 ;
  LAYER metal4 ;
  RECT 0.000 329.060 1.120 332.300 ;
  LAYER metal3 ;
  RECT 0.000 329.060 1.120 332.300 ;
  LAYER metal2 ;
  RECT 0.000 329.060 1.120 332.300 ;
  LAYER metal1 ;
  RECT 0.000 329.060 1.120 332.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 321.220 1.120 324.460 ;
  LAYER metal4 ;
  RECT 0.000 321.220 1.120 324.460 ;
  LAYER metal3 ;
  RECT 0.000 321.220 1.120 324.460 ;
  LAYER metal2 ;
  RECT 0.000 321.220 1.120 324.460 ;
  LAYER metal1 ;
  RECT 0.000 321.220 1.120 324.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 282.020 1.120 285.260 ;
  LAYER metal4 ;
  RECT 0.000 282.020 1.120 285.260 ;
  LAYER metal3 ;
  RECT 0.000 282.020 1.120 285.260 ;
  LAYER metal2 ;
  RECT 0.000 282.020 1.120 285.260 ;
  LAYER metal1 ;
  RECT 0.000 282.020 1.120 285.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 274.180 1.120 277.420 ;
  LAYER metal4 ;
  RECT 0.000 274.180 1.120 277.420 ;
  LAYER metal3 ;
  RECT 0.000 274.180 1.120 277.420 ;
  LAYER metal2 ;
  RECT 0.000 274.180 1.120 277.420 ;
  LAYER metal1 ;
  RECT 0.000 274.180 1.120 277.420 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 266.340 1.120 269.580 ;
  LAYER metal4 ;
  RECT 0.000 266.340 1.120 269.580 ;
  LAYER metal3 ;
  RECT 0.000 266.340 1.120 269.580 ;
  LAYER metal2 ;
  RECT 0.000 266.340 1.120 269.580 ;
  LAYER metal1 ;
  RECT 0.000 266.340 1.120 269.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 258.500 1.120 261.740 ;
  LAYER metal4 ;
  RECT 0.000 258.500 1.120 261.740 ;
  LAYER metal3 ;
  RECT 0.000 258.500 1.120 261.740 ;
  LAYER metal2 ;
  RECT 0.000 258.500 1.120 261.740 ;
  LAYER metal1 ;
  RECT 0.000 258.500 1.120 261.740 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 250.660 1.120 253.900 ;
  LAYER metal4 ;
  RECT 0.000 250.660 1.120 253.900 ;
  LAYER metal3 ;
  RECT 0.000 250.660 1.120 253.900 ;
  LAYER metal2 ;
  RECT 0.000 250.660 1.120 253.900 ;
  LAYER metal1 ;
  RECT 0.000 250.660 1.120 253.900 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 242.820 1.120 246.060 ;
  LAYER metal4 ;
  RECT 0.000 242.820 1.120 246.060 ;
  LAYER metal3 ;
  RECT 0.000 242.820 1.120 246.060 ;
  LAYER metal2 ;
  RECT 0.000 242.820 1.120 246.060 ;
  LAYER metal1 ;
  RECT 0.000 242.820 1.120 246.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 203.620 1.120 206.860 ;
  LAYER metal4 ;
  RECT 0.000 203.620 1.120 206.860 ;
  LAYER metal3 ;
  RECT 0.000 203.620 1.120 206.860 ;
  LAYER metal2 ;
  RECT 0.000 203.620 1.120 206.860 ;
  LAYER metal1 ;
  RECT 0.000 203.620 1.120 206.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 195.780 1.120 199.020 ;
  LAYER metal4 ;
  RECT 0.000 195.780 1.120 199.020 ;
  LAYER metal3 ;
  RECT 0.000 195.780 1.120 199.020 ;
  LAYER metal2 ;
  RECT 0.000 195.780 1.120 199.020 ;
  LAYER metal1 ;
  RECT 0.000 195.780 1.120 199.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 187.940 1.120 191.180 ;
  LAYER metal4 ;
  RECT 0.000 187.940 1.120 191.180 ;
  LAYER metal3 ;
  RECT 0.000 187.940 1.120 191.180 ;
  LAYER metal2 ;
  RECT 0.000 187.940 1.120 191.180 ;
  LAYER metal1 ;
  RECT 0.000 187.940 1.120 191.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 180.100 1.120 183.340 ;
  LAYER metal4 ;
  RECT 0.000 180.100 1.120 183.340 ;
  LAYER metal3 ;
  RECT 0.000 180.100 1.120 183.340 ;
  LAYER metal2 ;
  RECT 0.000 180.100 1.120 183.340 ;
  LAYER metal1 ;
  RECT 0.000 180.100 1.120 183.340 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 172.260 1.120 175.500 ;
  LAYER metal4 ;
  RECT 0.000 172.260 1.120 175.500 ;
  LAYER metal3 ;
  RECT 0.000 172.260 1.120 175.500 ;
  LAYER metal2 ;
  RECT 0.000 172.260 1.120 175.500 ;
  LAYER metal1 ;
  RECT 0.000 172.260 1.120 175.500 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 164.420 1.120 167.660 ;
  LAYER metal4 ;
  RECT 0.000 164.420 1.120 167.660 ;
  LAYER metal3 ;
  RECT 0.000 164.420 1.120 167.660 ;
  LAYER metal2 ;
  RECT 0.000 164.420 1.120 167.660 ;
  LAYER metal1 ;
  RECT 0.000 164.420 1.120 167.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 125.220 1.120 128.460 ;
  LAYER metal4 ;
  RECT 0.000 125.220 1.120 128.460 ;
  LAYER metal3 ;
  RECT 0.000 125.220 1.120 128.460 ;
  LAYER metal2 ;
  RECT 0.000 125.220 1.120 128.460 ;
  LAYER metal1 ;
  RECT 0.000 125.220 1.120 128.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 117.380 1.120 120.620 ;
  LAYER metal4 ;
  RECT 0.000 117.380 1.120 120.620 ;
  LAYER metal3 ;
  RECT 0.000 117.380 1.120 120.620 ;
  LAYER metal2 ;
  RECT 0.000 117.380 1.120 120.620 ;
  LAYER metal1 ;
  RECT 0.000 117.380 1.120 120.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 109.540 1.120 112.780 ;
  LAYER metal4 ;
  RECT 0.000 109.540 1.120 112.780 ;
  LAYER metal3 ;
  RECT 0.000 109.540 1.120 112.780 ;
  LAYER metal2 ;
  RECT 0.000 109.540 1.120 112.780 ;
  LAYER metal1 ;
  RECT 0.000 109.540 1.120 112.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 101.700 1.120 104.940 ;
  LAYER metal4 ;
  RECT 0.000 101.700 1.120 104.940 ;
  LAYER metal3 ;
  RECT 0.000 101.700 1.120 104.940 ;
  LAYER metal2 ;
  RECT 0.000 101.700 1.120 104.940 ;
  LAYER metal1 ;
  RECT 0.000 101.700 1.120 104.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 93.860 1.120 97.100 ;
  LAYER metal4 ;
  RECT 0.000 93.860 1.120 97.100 ;
  LAYER metal3 ;
  RECT 0.000 93.860 1.120 97.100 ;
  LAYER metal2 ;
  RECT 0.000 93.860 1.120 97.100 ;
  LAYER metal1 ;
  RECT 0.000 93.860 1.120 97.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 86.020 1.120 89.260 ;
  LAYER metal4 ;
  RECT 0.000 86.020 1.120 89.260 ;
  LAYER metal3 ;
  RECT 0.000 86.020 1.120 89.260 ;
  LAYER metal2 ;
  RECT 0.000 86.020 1.120 89.260 ;
  LAYER metal1 ;
  RECT 0.000 86.020 1.120 89.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 46.820 1.120 50.060 ;
  LAYER metal4 ;
  RECT 0.000 46.820 1.120 50.060 ;
  LAYER metal3 ;
  RECT 0.000 46.820 1.120 50.060 ;
  LAYER metal2 ;
  RECT 0.000 46.820 1.120 50.060 ;
  LAYER metal1 ;
  RECT 0.000 46.820 1.120 50.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 38.980 1.120 42.220 ;
  LAYER metal4 ;
  RECT 0.000 38.980 1.120 42.220 ;
  LAYER metal3 ;
  RECT 0.000 38.980 1.120 42.220 ;
  LAYER metal2 ;
  RECT 0.000 38.980 1.120 42.220 ;
  LAYER metal1 ;
  RECT 0.000 38.980 1.120 42.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 31.140 1.120 34.380 ;
  LAYER metal4 ;
  RECT 0.000 31.140 1.120 34.380 ;
  LAYER metal3 ;
  RECT 0.000 31.140 1.120 34.380 ;
  LAYER metal2 ;
  RECT 0.000 31.140 1.120 34.380 ;
  LAYER metal1 ;
  RECT 0.000 31.140 1.120 34.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 23.300 1.120 26.540 ;
  LAYER metal4 ;
  RECT 0.000 23.300 1.120 26.540 ;
  LAYER metal3 ;
  RECT 0.000 23.300 1.120 26.540 ;
  LAYER metal2 ;
  RECT 0.000 23.300 1.120 26.540 ;
  LAYER metal1 ;
  RECT 0.000 23.300 1.120 26.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 15.460 1.120 18.700 ;
  LAYER metal4 ;
  RECT 0.000 15.460 1.120 18.700 ;
  LAYER metal3 ;
  RECT 0.000 15.460 1.120 18.700 ;
  LAYER metal2 ;
  RECT 0.000 15.460 1.120 18.700 ;
  LAYER metal1 ;
  RECT 0.000 15.460 1.120 18.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 7.620 1.120 10.860 ;
  LAYER metal4 ;
  RECT 0.000 7.620 1.120 10.860 ;
  LAYER metal3 ;
  RECT 0.000 7.620 1.120 10.860 ;
  LAYER metal2 ;
  RECT 0.000 7.620 1.120 10.860 ;
  LAYER metal1 ;
  RECT 0.000 7.620 1.120 10.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3584.000 500.640 3587.540 501.760 ;
  LAYER metal4 ;
  RECT 3584.000 500.640 3587.540 501.760 ;
  LAYER metal3 ;
  RECT 3584.000 500.640 3587.540 501.760 ;
  LAYER metal2 ;
  RECT 3584.000 500.640 3587.540 501.760 ;
  LAYER metal1 ;
  RECT 3584.000 500.640 3587.540 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3575.320 500.640 3578.860 501.760 ;
  LAYER metal4 ;
  RECT 3575.320 500.640 3578.860 501.760 ;
  LAYER metal3 ;
  RECT 3575.320 500.640 3578.860 501.760 ;
  LAYER metal2 ;
  RECT 3575.320 500.640 3578.860 501.760 ;
  LAYER metal1 ;
  RECT 3575.320 500.640 3578.860 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3561.680 500.640 3565.220 501.760 ;
  LAYER metal4 ;
  RECT 3561.680 500.640 3565.220 501.760 ;
  LAYER metal3 ;
  RECT 3561.680 500.640 3565.220 501.760 ;
  LAYER metal2 ;
  RECT 3561.680 500.640 3565.220 501.760 ;
  LAYER metal1 ;
  RECT 3561.680 500.640 3565.220 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3548.660 500.640 3552.200 501.760 ;
  LAYER metal4 ;
  RECT 3548.660 500.640 3552.200 501.760 ;
  LAYER metal3 ;
  RECT 3548.660 500.640 3552.200 501.760 ;
  LAYER metal2 ;
  RECT 3548.660 500.640 3552.200 501.760 ;
  LAYER metal1 ;
  RECT 3548.660 500.640 3552.200 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3535.020 500.640 3538.560 501.760 ;
  LAYER metal4 ;
  RECT 3535.020 500.640 3538.560 501.760 ;
  LAYER metal3 ;
  RECT 3535.020 500.640 3538.560 501.760 ;
  LAYER metal2 ;
  RECT 3535.020 500.640 3538.560 501.760 ;
  LAYER metal1 ;
  RECT 3535.020 500.640 3538.560 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3521.380 500.640 3524.920 501.760 ;
  LAYER metal4 ;
  RECT 3521.380 500.640 3524.920 501.760 ;
  LAYER metal3 ;
  RECT 3521.380 500.640 3524.920 501.760 ;
  LAYER metal2 ;
  RECT 3521.380 500.640 3524.920 501.760 ;
  LAYER metal1 ;
  RECT 3521.380 500.640 3524.920 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3454.420 500.640 3457.960 501.760 ;
  LAYER metal4 ;
  RECT 3454.420 500.640 3457.960 501.760 ;
  LAYER metal3 ;
  RECT 3454.420 500.640 3457.960 501.760 ;
  LAYER metal2 ;
  RECT 3454.420 500.640 3457.960 501.760 ;
  LAYER metal1 ;
  RECT 3454.420 500.640 3457.960 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3440.780 500.640 3444.320 501.760 ;
  LAYER metal4 ;
  RECT 3440.780 500.640 3444.320 501.760 ;
  LAYER metal3 ;
  RECT 3440.780 500.640 3444.320 501.760 ;
  LAYER metal2 ;
  RECT 3440.780 500.640 3444.320 501.760 ;
  LAYER metal1 ;
  RECT 3440.780 500.640 3444.320 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3427.760 500.640 3431.300 501.760 ;
  LAYER metal4 ;
  RECT 3427.760 500.640 3431.300 501.760 ;
  LAYER metal3 ;
  RECT 3427.760 500.640 3431.300 501.760 ;
  LAYER metal2 ;
  RECT 3427.760 500.640 3431.300 501.760 ;
  LAYER metal1 ;
  RECT 3427.760 500.640 3431.300 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3414.120 500.640 3417.660 501.760 ;
  LAYER metal4 ;
  RECT 3414.120 500.640 3417.660 501.760 ;
  LAYER metal3 ;
  RECT 3414.120 500.640 3417.660 501.760 ;
  LAYER metal2 ;
  RECT 3414.120 500.640 3417.660 501.760 ;
  LAYER metal1 ;
  RECT 3414.120 500.640 3417.660 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3400.480 500.640 3404.020 501.760 ;
  LAYER metal4 ;
  RECT 3400.480 500.640 3404.020 501.760 ;
  LAYER metal3 ;
  RECT 3400.480 500.640 3404.020 501.760 ;
  LAYER metal2 ;
  RECT 3400.480 500.640 3404.020 501.760 ;
  LAYER metal1 ;
  RECT 3400.480 500.640 3404.020 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3387.460 500.640 3391.000 501.760 ;
  LAYER metal4 ;
  RECT 3387.460 500.640 3391.000 501.760 ;
  LAYER metal3 ;
  RECT 3387.460 500.640 3391.000 501.760 ;
  LAYER metal2 ;
  RECT 3387.460 500.640 3391.000 501.760 ;
  LAYER metal1 ;
  RECT 3387.460 500.640 3391.000 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3319.880 500.640 3323.420 501.760 ;
  LAYER metal4 ;
  RECT 3319.880 500.640 3323.420 501.760 ;
  LAYER metal3 ;
  RECT 3319.880 500.640 3323.420 501.760 ;
  LAYER metal2 ;
  RECT 3319.880 500.640 3323.420 501.760 ;
  LAYER metal1 ;
  RECT 3319.880 500.640 3323.420 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3306.860 500.640 3310.400 501.760 ;
  LAYER metal4 ;
  RECT 3306.860 500.640 3310.400 501.760 ;
  LAYER metal3 ;
  RECT 3306.860 500.640 3310.400 501.760 ;
  LAYER metal2 ;
  RECT 3306.860 500.640 3310.400 501.760 ;
  LAYER metal1 ;
  RECT 3306.860 500.640 3310.400 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3293.220 500.640 3296.760 501.760 ;
  LAYER metal4 ;
  RECT 3293.220 500.640 3296.760 501.760 ;
  LAYER metal3 ;
  RECT 3293.220 500.640 3296.760 501.760 ;
  LAYER metal2 ;
  RECT 3293.220 500.640 3296.760 501.760 ;
  LAYER metal1 ;
  RECT 3293.220 500.640 3296.760 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3279.580 500.640 3283.120 501.760 ;
  LAYER metal4 ;
  RECT 3279.580 500.640 3283.120 501.760 ;
  LAYER metal3 ;
  RECT 3279.580 500.640 3283.120 501.760 ;
  LAYER metal2 ;
  RECT 3279.580 500.640 3283.120 501.760 ;
  LAYER metal1 ;
  RECT 3279.580 500.640 3283.120 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3266.560 500.640 3270.100 501.760 ;
  LAYER metal4 ;
  RECT 3266.560 500.640 3270.100 501.760 ;
  LAYER metal3 ;
  RECT 3266.560 500.640 3270.100 501.760 ;
  LAYER metal2 ;
  RECT 3266.560 500.640 3270.100 501.760 ;
  LAYER metal1 ;
  RECT 3266.560 500.640 3270.100 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3252.920 500.640 3256.460 501.760 ;
  LAYER metal4 ;
  RECT 3252.920 500.640 3256.460 501.760 ;
  LAYER metal3 ;
  RECT 3252.920 500.640 3256.460 501.760 ;
  LAYER metal2 ;
  RECT 3252.920 500.640 3256.460 501.760 ;
  LAYER metal1 ;
  RECT 3252.920 500.640 3256.460 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3185.960 500.640 3189.500 501.760 ;
  LAYER metal4 ;
  RECT 3185.960 500.640 3189.500 501.760 ;
  LAYER metal3 ;
  RECT 3185.960 500.640 3189.500 501.760 ;
  LAYER metal2 ;
  RECT 3185.960 500.640 3189.500 501.760 ;
  LAYER metal1 ;
  RECT 3185.960 500.640 3189.500 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3172.320 500.640 3175.860 501.760 ;
  LAYER metal4 ;
  RECT 3172.320 500.640 3175.860 501.760 ;
  LAYER metal3 ;
  RECT 3172.320 500.640 3175.860 501.760 ;
  LAYER metal2 ;
  RECT 3172.320 500.640 3175.860 501.760 ;
  LAYER metal1 ;
  RECT 3172.320 500.640 3175.860 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3158.680 500.640 3162.220 501.760 ;
  LAYER metal4 ;
  RECT 3158.680 500.640 3162.220 501.760 ;
  LAYER metal3 ;
  RECT 3158.680 500.640 3162.220 501.760 ;
  LAYER metal2 ;
  RECT 3158.680 500.640 3162.220 501.760 ;
  LAYER metal1 ;
  RECT 3158.680 500.640 3162.220 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3145.040 500.640 3148.580 501.760 ;
  LAYER metal4 ;
  RECT 3145.040 500.640 3148.580 501.760 ;
  LAYER metal3 ;
  RECT 3145.040 500.640 3148.580 501.760 ;
  LAYER metal2 ;
  RECT 3145.040 500.640 3148.580 501.760 ;
  LAYER metal1 ;
  RECT 3145.040 500.640 3148.580 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3132.020 500.640 3135.560 501.760 ;
  LAYER metal4 ;
  RECT 3132.020 500.640 3135.560 501.760 ;
  LAYER metal3 ;
  RECT 3132.020 500.640 3135.560 501.760 ;
  LAYER metal2 ;
  RECT 3132.020 500.640 3135.560 501.760 ;
  LAYER metal1 ;
  RECT 3132.020 500.640 3135.560 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3118.380 500.640 3121.920 501.760 ;
  LAYER metal4 ;
  RECT 3118.380 500.640 3121.920 501.760 ;
  LAYER metal3 ;
  RECT 3118.380 500.640 3121.920 501.760 ;
  LAYER metal2 ;
  RECT 3118.380 500.640 3121.920 501.760 ;
  LAYER metal1 ;
  RECT 3118.380 500.640 3121.920 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3051.420 500.640 3054.960 501.760 ;
  LAYER metal4 ;
  RECT 3051.420 500.640 3054.960 501.760 ;
  LAYER metal3 ;
  RECT 3051.420 500.640 3054.960 501.760 ;
  LAYER metal2 ;
  RECT 3051.420 500.640 3054.960 501.760 ;
  LAYER metal1 ;
  RECT 3051.420 500.640 3054.960 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3037.780 500.640 3041.320 501.760 ;
  LAYER metal4 ;
  RECT 3037.780 500.640 3041.320 501.760 ;
  LAYER metal3 ;
  RECT 3037.780 500.640 3041.320 501.760 ;
  LAYER metal2 ;
  RECT 3037.780 500.640 3041.320 501.760 ;
  LAYER metal1 ;
  RECT 3037.780 500.640 3041.320 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3024.140 500.640 3027.680 501.760 ;
  LAYER metal4 ;
  RECT 3024.140 500.640 3027.680 501.760 ;
  LAYER metal3 ;
  RECT 3024.140 500.640 3027.680 501.760 ;
  LAYER metal2 ;
  RECT 3024.140 500.640 3027.680 501.760 ;
  LAYER metal1 ;
  RECT 3024.140 500.640 3027.680 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3011.120 500.640 3014.660 501.760 ;
  LAYER metal4 ;
  RECT 3011.120 500.640 3014.660 501.760 ;
  LAYER metal3 ;
  RECT 3011.120 500.640 3014.660 501.760 ;
  LAYER metal2 ;
  RECT 3011.120 500.640 3014.660 501.760 ;
  LAYER metal1 ;
  RECT 3011.120 500.640 3014.660 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2997.480 500.640 3001.020 501.760 ;
  LAYER metal4 ;
  RECT 2997.480 500.640 3001.020 501.760 ;
  LAYER metal3 ;
  RECT 2997.480 500.640 3001.020 501.760 ;
  LAYER metal2 ;
  RECT 2997.480 500.640 3001.020 501.760 ;
  LAYER metal1 ;
  RECT 2997.480 500.640 3001.020 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2983.840 500.640 2987.380 501.760 ;
  LAYER metal4 ;
  RECT 2983.840 500.640 2987.380 501.760 ;
  LAYER metal3 ;
  RECT 2983.840 500.640 2987.380 501.760 ;
  LAYER metal2 ;
  RECT 2983.840 500.640 2987.380 501.760 ;
  LAYER metal1 ;
  RECT 2983.840 500.640 2987.380 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2916.880 500.640 2920.420 501.760 ;
  LAYER metal4 ;
  RECT 2916.880 500.640 2920.420 501.760 ;
  LAYER metal3 ;
  RECT 2916.880 500.640 2920.420 501.760 ;
  LAYER metal2 ;
  RECT 2916.880 500.640 2920.420 501.760 ;
  LAYER metal1 ;
  RECT 2916.880 500.640 2920.420 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2903.240 500.640 2906.780 501.760 ;
  LAYER metal4 ;
  RECT 2903.240 500.640 2906.780 501.760 ;
  LAYER metal3 ;
  RECT 2903.240 500.640 2906.780 501.760 ;
  LAYER metal2 ;
  RECT 2903.240 500.640 2906.780 501.760 ;
  LAYER metal1 ;
  RECT 2903.240 500.640 2906.780 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2890.220 500.640 2893.760 501.760 ;
  LAYER metal4 ;
  RECT 2890.220 500.640 2893.760 501.760 ;
  LAYER metal3 ;
  RECT 2890.220 500.640 2893.760 501.760 ;
  LAYER metal2 ;
  RECT 2890.220 500.640 2893.760 501.760 ;
  LAYER metal1 ;
  RECT 2890.220 500.640 2893.760 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2876.580 500.640 2880.120 501.760 ;
  LAYER metal4 ;
  RECT 2876.580 500.640 2880.120 501.760 ;
  LAYER metal3 ;
  RECT 2876.580 500.640 2880.120 501.760 ;
  LAYER metal2 ;
  RECT 2876.580 500.640 2880.120 501.760 ;
  LAYER metal1 ;
  RECT 2876.580 500.640 2880.120 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2862.940 500.640 2866.480 501.760 ;
  LAYER metal4 ;
  RECT 2862.940 500.640 2866.480 501.760 ;
  LAYER metal3 ;
  RECT 2862.940 500.640 2866.480 501.760 ;
  LAYER metal2 ;
  RECT 2862.940 500.640 2866.480 501.760 ;
  LAYER metal1 ;
  RECT 2862.940 500.640 2866.480 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2849.920 500.640 2853.460 501.760 ;
  LAYER metal4 ;
  RECT 2849.920 500.640 2853.460 501.760 ;
  LAYER metal3 ;
  RECT 2849.920 500.640 2853.460 501.760 ;
  LAYER metal2 ;
  RECT 2849.920 500.640 2853.460 501.760 ;
  LAYER metal1 ;
  RECT 2849.920 500.640 2853.460 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2782.340 500.640 2785.880 501.760 ;
  LAYER metal4 ;
  RECT 2782.340 500.640 2785.880 501.760 ;
  LAYER metal3 ;
  RECT 2782.340 500.640 2785.880 501.760 ;
  LAYER metal2 ;
  RECT 2782.340 500.640 2785.880 501.760 ;
  LAYER metal1 ;
  RECT 2782.340 500.640 2785.880 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2769.320 500.640 2772.860 501.760 ;
  LAYER metal4 ;
  RECT 2769.320 500.640 2772.860 501.760 ;
  LAYER metal3 ;
  RECT 2769.320 500.640 2772.860 501.760 ;
  LAYER metal2 ;
  RECT 2769.320 500.640 2772.860 501.760 ;
  LAYER metal1 ;
  RECT 2769.320 500.640 2772.860 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2755.680 500.640 2759.220 501.760 ;
  LAYER metal4 ;
  RECT 2755.680 500.640 2759.220 501.760 ;
  LAYER metal3 ;
  RECT 2755.680 500.640 2759.220 501.760 ;
  LAYER metal2 ;
  RECT 2755.680 500.640 2759.220 501.760 ;
  LAYER metal1 ;
  RECT 2755.680 500.640 2759.220 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2742.040 500.640 2745.580 501.760 ;
  LAYER metal4 ;
  RECT 2742.040 500.640 2745.580 501.760 ;
  LAYER metal3 ;
  RECT 2742.040 500.640 2745.580 501.760 ;
  LAYER metal2 ;
  RECT 2742.040 500.640 2745.580 501.760 ;
  LAYER metal1 ;
  RECT 2742.040 500.640 2745.580 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2728.400 500.640 2731.940 501.760 ;
  LAYER metal4 ;
  RECT 2728.400 500.640 2731.940 501.760 ;
  LAYER metal3 ;
  RECT 2728.400 500.640 2731.940 501.760 ;
  LAYER metal2 ;
  RECT 2728.400 500.640 2731.940 501.760 ;
  LAYER metal1 ;
  RECT 2728.400 500.640 2731.940 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2715.380 500.640 2718.920 501.760 ;
  LAYER metal4 ;
  RECT 2715.380 500.640 2718.920 501.760 ;
  LAYER metal3 ;
  RECT 2715.380 500.640 2718.920 501.760 ;
  LAYER metal2 ;
  RECT 2715.380 500.640 2718.920 501.760 ;
  LAYER metal1 ;
  RECT 2715.380 500.640 2718.920 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2647.800 500.640 2651.340 501.760 ;
  LAYER metal4 ;
  RECT 2647.800 500.640 2651.340 501.760 ;
  LAYER metal3 ;
  RECT 2647.800 500.640 2651.340 501.760 ;
  LAYER metal2 ;
  RECT 2647.800 500.640 2651.340 501.760 ;
  LAYER metal1 ;
  RECT 2647.800 500.640 2651.340 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2634.780 500.640 2638.320 501.760 ;
  LAYER metal4 ;
  RECT 2634.780 500.640 2638.320 501.760 ;
  LAYER metal3 ;
  RECT 2634.780 500.640 2638.320 501.760 ;
  LAYER metal2 ;
  RECT 2634.780 500.640 2638.320 501.760 ;
  LAYER metal1 ;
  RECT 2634.780 500.640 2638.320 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2621.140 500.640 2624.680 501.760 ;
  LAYER metal4 ;
  RECT 2621.140 500.640 2624.680 501.760 ;
  LAYER metal3 ;
  RECT 2621.140 500.640 2624.680 501.760 ;
  LAYER metal2 ;
  RECT 2621.140 500.640 2624.680 501.760 ;
  LAYER metal1 ;
  RECT 2621.140 500.640 2624.680 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2607.500 500.640 2611.040 501.760 ;
  LAYER metal4 ;
  RECT 2607.500 500.640 2611.040 501.760 ;
  LAYER metal3 ;
  RECT 2607.500 500.640 2611.040 501.760 ;
  LAYER metal2 ;
  RECT 2607.500 500.640 2611.040 501.760 ;
  LAYER metal1 ;
  RECT 2607.500 500.640 2611.040 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2594.480 500.640 2598.020 501.760 ;
  LAYER metal4 ;
  RECT 2594.480 500.640 2598.020 501.760 ;
  LAYER metal3 ;
  RECT 2594.480 500.640 2598.020 501.760 ;
  LAYER metal2 ;
  RECT 2594.480 500.640 2598.020 501.760 ;
  LAYER metal1 ;
  RECT 2594.480 500.640 2598.020 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2580.840 500.640 2584.380 501.760 ;
  LAYER metal4 ;
  RECT 2580.840 500.640 2584.380 501.760 ;
  LAYER metal3 ;
  RECT 2580.840 500.640 2584.380 501.760 ;
  LAYER metal2 ;
  RECT 2580.840 500.640 2584.380 501.760 ;
  LAYER metal1 ;
  RECT 2580.840 500.640 2584.380 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2513.880 500.640 2517.420 501.760 ;
  LAYER metal4 ;
  RECT 2513.880 500.640 2517.420 501.760 ;
  LAYER metal3 ;
  RECT 2513.880 500.640 2517.420 501.760 ;
  LAYER metal2 ;
  RECT 2513.880 500.640 2517.420 501.760 ;
  LAYER metal1 ;
  RECT 2513.880 500.640 2517.420 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2500.240 500.640 2503.780 501.760 ;
  LAYER metal4 ;
  RECT 2500.240 500.640 2503.780 501.760 ;
  LAYER metal3 ;
  RECT 2500.240 500.640 2503.780 501.760 ;
  LAYER metal2 ;
  RECT 2500.240 500.640 2503.780 501.760 ;
  LAYER metal1 ;
  RECT 2500.240 500.640 2503.780 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2486.600 500.640 2490.140 501.760 ;
  LAYER metal4 ;
  RECT 2486.600 500.640 2490.140 501.760 ;
  LAYER metal3 ;
  RECT 2486.600 500.640 2490.140 501.760 ;
  LAYER metal2 ;
  RECT 2486.600 500.640 2490.140 501.760 ;
  LAYER metal1 ;
  RECT 2486.600 500.640 2490.140 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2473.580 500.640 2477.120 501.760 ;
  LAYER metal4 ;
  RECT 2473.580 500.640 2477.120 501.760 ;
  LAYER metal3 ;
  RECT 2473.580 500.640 2477.120 501.760 ;
  LAYER metal2 ;
  RECT 2473.580 500.640 2477.120 501.760 ;
  LAYER metal1 ;
  RECT 2473.580 500.640 2477.120 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2459.940 500.640 2463.480 501.760 ;
  LAYER metal4 ;
  RECT 2459.940 500.640 2463.480 501.760 ;
  LAYER metal3 ;
  RECT 2459.940 500.640 2463.480 501.760 ;
  LAYER metal2 ;
  RECT 2459.940 500.640 2463.480 501.760 ;
  LAYER metal1 ;
  RECT 2459.940 500.640 2463.480 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2446.300 500.640 2449.840 501.760 ;
  LAYER metal4 ;
  RECT 2446.300 500.640 2449.840 501.760 ;
  LAYER metal3 ;
  RECT 2446.300 500.640 2449.840 501.760 ;
  LAYER metal2 ;
  RECT 2446.300 500.640 2449.840 501.760 ;
  LAYER metal1 ;
  RECT 2446.300 500.640 2449.840 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2379.340 500.640 2382.880 501.760 ;
  LAYER metal4 ;
  RECT 2379.340 500.640 2382.880 501.760 ;
  LAYER metal3 ;
  RECT 2379.340 500.640 2382.880 501.760 ;
  LAYER metal2 ;
  RECT 2379.340 500.640 2382.880 501.760 ;
  LAYER metal1 ;
  RECT 2379.340 500.640 2382.880 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2365.700 500.640 2369.240 501.760 ;
  LAYER metal4 ;
  RECT 2365.700 500.640 2369.240 501.760 ;
  LAYER metal3 ;
  RECT 2365.700 500.640 2369.240 501.760 ;
  LAYER metal2 ;
  RECT 2365.700 500.640 2369.240 501.760 ;
  LAYER metal1 ;
  RECT 2365.700 500.640 2369.240 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2352.680 500.640 2356.220 501.760 ;
  LAYER metal4 ;
  RECT 2352.680 500.640 2356.220 501.760 ;
  LAYER metal3 ;
  RECT 2352.680 500.640 2356.220 501.760 ;
  LAYER metal2 ;
  RECT 2352.680 500.640 2356.220 501.760 ;
  LAYER metal1 ;
  RECT 2352.680 500.640 2356.220 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2339.040 500.640 2342.580 501.760 ;
  LAYER metal4 ;
  RECT 2339.040 500.640 2342.580 501.760 ;
  LAYER metal3 ;
  RECT 2339.040 500.640 2342.580 501.760 ;
  LAYER metal2 ;
  RECT 2339.040 500.640 2342.580 501.760 ;
  LAYER metal1 ;
  RECT 2339.040 500.640 2342.580 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2325.400 500.640 2328.940 501.760 ;
  LAYER metal4 ;
  RECT 2325.400 500.640 2328.940 501.760 ;
  LAYER metal3 ;
  RECT 2325.400 500.640 2328.940 501.760 ;
  LAYER metal2 ;
  RECT 2325.400 500.640 2328.940 501.760 ;
  LAYER metal1 ;
  RECT 2325.400 500.640 2328.940 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2311.760 500.640 2315.300 501.760 ;
  LAYER metal4 ;
  RECT 2311.760 500.640 2315.300 501.760 ;
  LAYER metal3 ;
  RECT 2311.760 500.640 2315.300 501.760 ;
  LAYER metal2 ;
  RECT 2311.760 500.640 2315.300 501.760 ;
  LAYER metal1 ;
  RECT 2311.760 500.640 2315.300 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2244.800 500.640 2248.340 501.760 ;
  LAYER metal4 ;
  RECT 2244.800 500.640 2248.340 501.760 ;
  LAYER metal3 ;
  RECT 2244.800 500.640 2248.340 501.760 ;
  LAYER metal2 ;
  RECT 2244.800 500.640 2248.340 501.760 ;
  LAYER metal1 ;
  RECT 2244.800 500.640 2248.340 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2231.160 500.640 2234.700 501.760 ;
  LAYER metal4 ;
  RECT 2231.160 500.640 2234.700 501.760 ;
  LAYER metal3 ;
  RECT 2231.160 500.640 2234.700 501.760 ;
  LAYER metal2 ;
  RECT 2231.160 500.640 2234.700 501.760 ;
  LAYER metal1 ;
  RECT 2231.160 500.640 2234.700 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2218.140 500.640 2221.680 501.760 ;
  LAYER metal4 ;
  RECT 2218.140 500.640 2221.680 501.760 ;
  LAYER metal3 ;
  RECT 2218.140 500.640 2221.680 501.760 ;
  LAYER metal2 ;
  RECT 2218.140 500.640 2221.680 501.760 ;
  LAYER metal1 ;
  RECT 2218.140 500.640 2221.680 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2204.500 500.640 2208.040 501.760 ;
  LAYER metal4 ;
  RECT 2204.500 500.640 2208.040 501.760 ;
  LAYER metal3 ;
  RECT 2204.500 500.640 2208.040 501.760 ;
  LAYER metal2 ;
  RECT 2204.500 500.640 2208.040 501.760 ;
  LAYER metal1 ;
  RECT 2204.500 500.640 2208.040 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2190.860 500.640 2194.400 501.760 ;
  LAYER metal4 ;
  RECT 2190.860 500.640 2194.400 501.760 ;
  LAYER metal3 ;
  RECT 2190.860 500.640 2194.400 501.760 ;
  LAYER metal2 ;
  RECT 2190.860 500.640 2194.400 501.760 ;
  LAYER metal1 ;
  RECT 2190.860 500.640 2194.400 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2177.840 500.640 2181.380 501.760 ;
  LAYER metal4 ;
  RECT 2177.840 500.640 2181.380 501.760 ;
  LAYER metal3 ;
  RECT 2177.840 500.640 2181.380 501.760 ;
  LAYER metal2 ;
  RECT 2177.840 500.640 2181.380 501.760 ;
  LAYER metal1 ;
  RECT 2177.840 500.640 2181.380 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2110.260 500.640 2113.800 501.760 ;
  LAYER metal4 ;
  RECT 2110.260 500.640 2113.800 501.760 ;
  LAYER metal3 ;
  RECT 2110.260 500.640 2113.800 501.760 ;
  LAYER metal2 ;
  RECT 2110.260 500.640 2113.800 501.760 ;
  LAYER metal1 ;
  RECT 2110.260 500.640 2113.800 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2097.240 500.640 2100.780 501.760 ;
  LAYER metal4 ;
  RECT 2097.240 500.640 2100.780 501.760 ;
  LAYER metal3 ;
  RECT 2097.240 500.640 2100.780 501.760 ;
  LAYER metal2 ;
  RECT 2097.240 500.640 2100.780 501.760 ;
  LAYER metal1 ;
  RECT 2097.240 500.640 2100.780 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2083.600 500.640 2087.140 501.760 ;
  LAYER metal4 ;
  RECT 2083.600 500.640 2087.140 501.760 ;
  LAYER metal3 ;
  RECT 2083.600 500.640 2087.140 501.760 ;
  LAYER metal2 ;
  RECT 2083.600 500.640 2087.140 501.760 ;
  LAYER metal1 ;
  RECT 2083.600 500.640 2087.140 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2069.960 500.640 2073.500 501.760 ;
  LAYER metal4 ;
  RECT 2069.960 500.640 2073.500 501.760 ;
  LAYER metal3 ;
  RECT 2069.960 500.640 2073.500 501.760 ;
  LAYER metal2 ;
  RECT 2069.960 500.640 2073.500 501.760 ;
  LAYER metal1 ;
  RECT 2069.960 500.640 2073.500 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2056.940 500.640 2060.480 501.760 ;
  LAYER metal4 ;
  RECT 2056.940 500.640 2060.480 501.760 ;
  LAYER metal3 ;
  RECT 2056.940 500.640 2060.480 501.760 ;
  LAYER metal2 ;
  RECT 2056.940 500.640 2060.480 501.760 ;
  LAYER metal1 ;
  RECT 2056.940 500.640 2060.480 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2043.300 500.640 2046.840 501.760 ;
  LAYER metal4 ;
  RECT 2043.300 500.640 2046.840 501.760 ;
  LAYER metal3 ;
  RECT 2043.300 500.640 2046.840 501.760 ;
  LAYER metal2 ;
  RECT 2043.300 500.640 2046.840 501.760 ;
  LAYER metal1 ;
  RECT 2043.300 500.640 2046.840 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1976.340 500.640 1979.880 501.760 ;
  LAYER metal4 ;
  RECT 1976.340 500.640 1979.880 501.760 ;
  LAYER metal3 ;
  RECT 1976.340 500.640 1979.880 501.760 ;
  LAYER metal2 ;
  RECT 1976.340 500.640 1979.880 501.760 ;
  LAYER metal1 ;
  RECT 1976.340 500.640 1979.880 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1962.700 500.640 1966.240 501.760 ;
  LAYER metal4 ;
  RECT 1962.700 500.640 1966.240 501.760 ;
  LAYER metal3 ;
  RECT 1962.700 500.640 1966.240 501.760 ;
  LAYER metal2 ;
  RECT 1962.700 500.640 1966.240 501.760 ;
  LAYER metal1 ;
  RECT 1962.700 500.640 1966.240 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1949.060 500.640 1952.600 501.760 ;
  LAYER metal4 ;
  RECT 1949.060 500.640 1952.600 501.760 ;
  LAYER metal3 ;
  RECT 1949.060 500.640 1952.600 501.760 ;
  LAYER metal2 ;
  RECT 1949.060 500.640 1952.600 501.760 ;
  LAYER metal1 ;
  RECT 1949.060 500.640 1952.600 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1936.040 500.640 1939.580 501.760 ;
  LAYER metal4 ;
  RECT 1936.040 500.640 1939.580 501.760 ;
  LAYER metal3 ;
  RECT 1936.040 500.640 1939.580 501.760 ;
  LAYER metal2 ;
  RECT 1936.040 500.640 1939.580 501.760 ;
  LAYER metal1 ;
  RECT 1936.040 500.640 1939.580 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1922.400 500.640 1925.940 501.760 ;
  LAYER metal4 ;
  RECT 1922.400 500.640 1925.940 501.760 ;
  LAYER metal3 ;
  RECT 1922.400 500.640 1925.940 501.760 ;
  LAYER metal2 ;
  RECT 1922.400 500.640 1925.940 501.760 ;
  LAYER metal1 ;
  RECT 1922.400 500.640 1925.940 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1908.760 500.640 1912.300 501.760 ;
  LAYER metal4 ;
  RECT 1908.760 500.640 1912.300 501.760 ;
  LAYER metal3 ;
  RECT 1908.760 500.640 1912.300 501.760 ;
  LAYER metal2 ;
  RECT 1908.760 500.640 1912.300 501.760 ;
  LAYER metal1 ;
  RECT 1908.760 500.640 1912.300 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1846.140 500.640 1849.680 501.760 ;
  LAYER metal4 ;
  RECT 1846.140 500.640 1849.680 501.760 ;
  LAYER metal3 ;
  RECT 1846.140 500.640 1849.680 501.760 ;
  LAYER metal2 ;
  RECT 1846.140 500.640 1849.680 501.760 ;
  LAYER metal1 ;
  RECT 1846.140 500.640 1849.680 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1833.120 500.640 1836.660 501.760 ;
  LAYER metal4 ;
  RECT 1833.120 500.640 1836.660 501.760 ;
  LAYER metal3 ;
  RECT 1833.120 500.640 1836.660 501.760 ;
  LAYER metal2 ;
  RECT 1833.120 500.640 1836.660 501.760 ;
  LAYER metal1 ;
  RECT 1833.120 500.640 1836.660 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1803.980 500.640 1807.520 501.760 ;
  LAYER metal4 ;
  RECT 1803.980 500.640 1807.520 501.760 ;
  LAYER metal3 ;
  RECT 1803.980 500.640 1807.520 501.760 ;
  LAYER metal2 ;
  RECT 1803.980 500.640 1807.520 501.760 ;
  LAYER metal1 ;
  RECT 1803.980 500.640 1807.520 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1779.800 500.640 1783.340 501.760 ;
  LAYER metal4 ;
  RECT 1779.800 500.640 1783.340 501.760 ;
  LAYER metal3 ;
  RECT 1779.800 500.640 1783.340 501.760 ;
  LAYER metal2 ;
  RECT 1779.800 500.640 1783.340 501.760 ;
  LAYER metal1 ;
  RECT 1779.800 500.640 1783.340 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1756.860 500.640 1760.400 501.760 ;
  LAYER metal4 ;
  RECT 1756.860 500.640 1760.400 501.760 ;
  LAYER metal3 ;
  RECT 1756.860 500.640 1760.400 501.760 ;
  LAYER metal2 ;
  RECT 1756.860 500.640 1760.400 501.760 ;
  LAYER metal1 ;
  RECT 1756.860 500.640 1760.400 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1748.180 500.640 1751.720 501.760 ;
  LAYER metal4 ;
  RECT 1748.180 500.640 1751.720 501.760 ;
  LAYER metal3 ;
  RECT 1748.180 500.640 1751.720 501.760 ;
  LAYER metal2 ;
  RECT 1748.180 500.640 1751.720 501.760 ;
  LAYER metal1 ;
  RECT 1748.180 500.640 1751.720 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1685.560 500.640 1689.100 501.760 ;
  LAYER metal4 ;
  RECT 1685.560 500.640 1689.100 501.760 ;
  LAYER metal3 ;
  RECT 1685.560 500.640 1689.100 501.760 ;
  LAYER metal2 ;
  RECT 1685.560 500.640 1689.100 501.760 ;
  LAYER metal1 ;
  RECT 1685.560 500.640 1689.100 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1672.540 500.640 1676.080 501.760 ;
  LAYER metal4 ;
  RECT 1672.540 500.640 1676.080 501.760 ;
  LAYER metal3 ;
  RECT 1672.540 500.640 1676.080 501.760 ;
  LAYER metal2 ;
  RECT 1672.540 500.640 1676.080 501.760 ;
  LAYER metal1 ;
  RECT 1672.540 500.640 1676.080 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1658.900 500.640 1662.440 501.760 ;
  LAYER metal4 ;
  RECT 1658.900 500.640 1662.440 501.760 ;
  LAYER metal3 ;
  RECT 1658.900 500.640 1662.440 501.760 ;
  LAYER metal2 ;
  RECT 1658.900 500.640 1662.440 501.760 ;
  LAYER metal1 ;
  RECT 1658.900 500.640 1662.440 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1645.260 500.640 1648.800 501.760 ;
  LAYER metal4 ;
  RECT 1645.260 500.640 1648.800 501.760 ;
  LAYER metal3 ;
  RECT 1645.260 500.640 1648.800 501.760 ;
  LAYER metal2 ;
  RECT 1645.260 500.640 1648.800 501.760 ;
  LAYER metal1 ;
  RECT 1645.260 500.640 1648.800 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1632.240 500.640 1635.780 501.760 ;
  LAYER metal4 ;
  RECT 1632.240 500.640 1635.780 501.760 ;
  LAYER metal3 ;
  RECT 1632.240 500.640 1635.780 501.760 ;
  LAYER metal2 ;
  RECT 1632.240 500.640 1635.780 501.760 ;
  LAYER metal1 ;
  RECT 1632.240 500.640 1635.780 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1618.600 500.640 1622.140 501.760 ;
  LAYER metal4 ;
  RECT 1618.600 500.640 1622.140 501.760 ;
  LAYER metal3 ;
  RECT 1618.600 500.640 1622.140 501.760 ;
  LAYER metal2 ;
  RECT 1618.600 500.640 1622.140 501.760 ;
  LAYER metal1 ;
  RECT 1618.600 500.640 1622.140 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1551.640 500.640 1555.180 501.760 ;
  LAYER metal4 ;
  RECT 1551.640 500.640 1555.180 501.760 ;
  LAYER metal3 ;
  RECT 1551.640 500.640 1555.180 501.760 ;
  LAYER metal2 ;
  RECT 1551.640 500.640 1555.180 501.760 ;
  LAYER metal1 ;
  RECT 1551.640 500.640 1555.180 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1538.000 500.640 1541.540 501.760 ;
  LAYER metal4 ;
  RECT 1538.000 500.640 1541.540 501.760 ;
  LAYER metal3 ;
  RECT 1538.000 500.640 1541.540 501.760 ;
  LAYER metal2 ;
  RECT 1538.000 500.640 1541.540 501.760 ;
  LAYER metal1 ;
  RECT 1538.000 500.640 1541.540 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1524.360 500.640 1527.900 501.760 ;
  LAYER metal4 ;
  RECT 1524.360 500.640 1527.900 501.760 ;
  LAYER metal3 ;
  RECT 1524.360 500.640 1527.900 501.760 ;
  LAYER metal2 ;
  RECT 1524.360 500.640 1527.900 501.760 ;
  LAYER metal1 ;
  RECT 1524.360 500.640 1527.900 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1511.340 500.640 1514.880 501.760 ;
  LAYER metal4 ;
  RECT 1511.340 500.640 1514.880 501.760 ;
  LAYER metal3 ;
  RECT 1511.340 500.640 1514.880 501.760 ;
  LAYER metal2 ;
  RECT 1511.340 500.640 1514.880 501.760 ;
  LAYER metal1 ;
  RECT 1511.340 500.640 1514.880 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1497.700 500.640 1501.240 501.760 ;
  LAYER metal4 ;
  RECT 1497.700 500.640 1501.240 501.760 ;
  LAYER metal3 ;
  RECT 1497.700 500.640 1501.240 501.760 ;
  LAYER metal2 ;
  RECT 1497.700 500.640 1501.240 501.760 ;
  LAYER metal1 ;
  RECT 1497.700 500.640 1501.240 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1484.060 500.640 1487.600 501.760 ;
  LAYER metal4 ;
  RECT 1484.060 500.640 1487.600 501.760 ;
  LAYER metal3 ;
  RECT 1484.060 500.640 1487.600 501.760 ;
  LAYER metal2 ;
  RECT 1484.060 500.640 1487.600 501.760 ;
  LAYER metal1 ;
  RECT 1484.060 500.640 1487.600 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1417.100 500.640 1420.640 501.760 ;
  LAYER metal4 ;
  RECT 1417.100 500.640 1420.640 501.760 ;
  LAYER metal3 ;
  RECT 1417.100 500.640 1420.640 501.760 ;
  LAYER metal2 ;
  RECT 1417.100 500.640 1420.640 501.760 ;
  LAYER metal1 ;
  RECT 1417.100 500.640 1420.640 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1403.460 500.640 1407.000 501.760 ;
  LAYER metal4 ;
  RECT 1403.460 500.640 1407.000 501.760 ;
  LAYER metal3 ;
  RECT 1403.460 500.640 1407.000 501.760 ;
  LAYER metal2 ;
  RECT 1403.460 500.640 1407.000 501.760 ;
  LAYER metal1 ;
  RECT 1403.460 500.640 1407.000 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1390.440 500.640 1393.980 501.760 ;
  LAYER metal4 ;
  RECT 1390.440 500.640 1393.980 501.760 ;
  LAYER metal3 ;
  RECT 1390.440 500.640 1393.980 501.760 ;
  LAYER metal2 ;
  RECT 1390.440 500.640 1393.980 501.760 ;
  LAYER metal1 ;
  RECT 1390.440 500.640 1393.980 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1376.800 500.640 1380.340 501.760 ;
  LAYER metal4 ;
  RECT 1376.800 500.640 1380.340 501.760 ;
  LAYER metal3 ;
  RECT 1376.800 500.640 1380.340 501.760 ;
  LAYER metal2 ;
  RECT 1376.800 500.640 1380.340 501.760 ;
  LAYER metal1 ;
  RECT 1376.800 500.640 1380.340 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1363.160 500.640 1366.700 501.760 ;
  LAYER metal4 ;
  RECT 1363.160 500.640 1366.700 501.760 ;
  LAYER metal3 ;
  RECT 1363.160 500.640 1366.700 501.760 ;
  LAYER metal2 ;
  RECT 1363.160 500.640 1366.700 501.760 ;
  LAYER metal1 ;
  RECT 1363.160 500.640 1366.700 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1350.140 500.640 1353.680 501.760 ;
  LAYER metal4 ;
  RECT 1350.140 500.640 1353.680 501.760 ;
  LAYER metal3 ;
  RECT 1350.140 500.640 1353.680 501.760 ;
  LAYER metal2 ;
  RECT 1350.140 500.640 1353.680 501.760 ;
  LAYER metal1 ;
  RECT 1350.140 500.640 1353.680 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1282.560 500.640 1286.100 501.760 ;
  LAYER metal4 ;
  RECT 1282.560 500.640 1286.100 501.760 ;
  LAYER metal3 ;
  RECT 1282.560 500.640 1286.100 501.760 ;
  LAYER metal2 ;
  RECT 1282.560 500.640 1286.100 501.760 ;
  LAYER metal1 ;
  RECT 1282.560 500.640 1286.100 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1268.920 500.640 1272.460 501.760 ;
  LAYER metal4 ;
  RECT 1268.920 500.640 1272.460 501.760 ;
  LAYER metal3 ;
  RECT 1268.920 500.640 1272.460 501.760 ;
  LAYER metal2 ;
  RECT 1268.920 500.640 1272.460 501.760 ;
  LAYER metal1 ;
  RECT 1268.920 500.640 1272.460 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1255.900 500.640 1259.440 501.760 ;
  LAYER metal4 ;
  RECT 1255.900 500.640 1259.440 501.760 ;
  LAYER metal3 ;
  RECT 1255.900 500.640 1259.440 501.760 ;
  LAYER metal2 ;
  RECT 1255.900 500.640 1259.440 501.760 ;
  LAYER metal1 ;
  RECT 1255.900 500.640 1259.440 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1242.260 500.640 1245.800 501.760 ;
  LAYER metal4 ;
  RECT 1242.260 500.640 1245.800 501.760 ;
  LAYER metal3 ;
  RECT 1242.260 500.640 1245.800 501.760 ;
  LAYER metal2 ;
  RECT 1242.260 500.640 1245.800 501.760 ;
  LAYER metal1 ;
  RECT 1242.260 500.640 1245.800 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1228.620 500.640 1232.160 501.760 ;
  LAYER metal4 ;
  RECT 1228.620 500.640 1232.160 501.760 ;
  LAYER metal3 ;
  RECT 1228.620 500.640 1232.160 501.760 ;
  LAYER metal2 ;
  RECT 1228.620 500.640 1232.160 501.760 ;
  LAYER metal1 ;
  RECT 1228.620 500.640 1232.160 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1215.600 500.640 1219.140 501.760 ;
  LAYER metal4 ;
  RECT 1215.600 500.640 1219.140 501.760 ;
  LAYER metal3 ;
  RECT 1215.600 500.640 1219.140 501.760 ;
  LAYER metal2 ;
  RECT 1215.600 500.640 1219.140 501.760 ;
  LAYER metal1 ;
  RECT 1215.600 500.640 1219.140 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1148.020 500.640 1151.560 501.760 ;
  LAYER metal4 ;
  RECT 1148.020 500.640 1151.560 501.760 ;
  LAYER metal3 ;
  RECT 1148.020 500.640 1151.560 501.760 ;
  LAYER metal2 ;
  RECT 1148.020 500.640 1151.560 501.760 ;
  LAYER metal1 ;
  RECT 1148.020 500.640 1151.560 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1135.000 500.640 1138.540 501.760 ;
  LAYER metal4 ;
  RECT 1135.000 500.640 1138.540 501.760 ;
  LAYER metal3 ;
  RECT 1135.000 500.640 1138.540 501.760 ;
  LAYER metal2 ;
  RECT 1135.000 500.640 1138.540 501.760 ;
  LAYER metal1 ;
  RECT 1135.000 500.640 1138.540 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1121.360 500.640 1124.900 501.760 ;
  LAYER metal4 ;
  RECT 1121.360 500.640 1124.900 501.760 ;
  LAYER metal3 ;
  RECT 1121.360 500.640 1124.900 501.760 ;
  LAYER metal2 ;
  RECT 1121.360 500.640 1124.900 501.760 ;
  LAYER metal1 ;
  RECT 1121.360 500.640 1124.900 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1107.720 500.640 1111.260 501.760 ;
  LAYER metal4 ;
  RECT 1107.720 500.640 1111.260 501.760 ;
  LAYER metal3 ;
  RECT 1107.720 500.640 1111.260 501.760 ;
  LAYER metal2 ;
  RECT 1107.720 500.640 1111.260 501.760 ;
  LAYER metal1 ;
  RECT 1107.720 500.640 1111.260 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1094.700 500.640 1098.240 501.760 ;
  LAYER metal4 ;
  RECT 1094.700 500.640 1098.240 501.760 ;
  LAYER metal3 ;
  RECT 1094.700 500.640 1098.240 501.760 ;
  LAYER metal2 ;
  RECT 1094.700 500.640 1098.240 501.760 ;
  LAYER metal1 ;
  RECT 1094.700 500.640 1098.240 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1081.060 500.640 1084.600 501.760 ;
  LAYER metal4 ;
  RECT 1081.060 500.640 1084.600 501.760 ;
  LAYER metal3 ;
  RECT 1081.060 500.640 1084.600 501.760 ;
  LAYER metal2 ;
  RECT 1081.060 500.640 1084.600 501.760 ;
  LAYER metal1 ;
  RECT 1081.060 500.640 1084.600 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1014.100 500.640 1017.640 501.760 ;
  LAYER metal4 ;
  RECT 1014.100 500.640 1017.640 501.760 ;
  LAYER metal3 ;
  RECT 1014.100 500.640 1017.640 501.760 ;
  LAYER metal2 ;
  RECT 1014.100 500.640 1017.640 501.760 ;
  LAYER metal1 ;
  RECT 1014.100 500.640 1017.640 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1000.460 500.640 1004.000 501.760 ;
  LAYER metal4 ;
  RECT 1000.460 500.640 1004.000 501.760 ;
  LAYER metal3 ;
  RECT 1000.460 500.640 1004.000 501.760 ;
  LAYER metal2 ;
  RECT 1000.460 500.640 1004.000 501.760 ;
  LAYER metal1 ;
  RECT 1000.460 500.640 1004.000 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 986.820 500.640 990.360 501.760 ;
  LAYER metal4 ;
  RECT 986.820 500.640 990.360 501.760 ;
  LAYER metal3 ;
  RECT 986.820 500.640 990.360 501.760 ;
  LAYER metal2 ;
  RECT 986.820 500.640 990.360 501.760 ;
  LAYER metal1 ;
  RECT 986.820 500.640 990.360 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 973.800 500.640 977.340 501.760 ;
  LAYER metal4 ;
  RECT 973.800 500.640 977.340 501.760 ;
  LAYER metal3 ;
  RECT 973.800 500.640 977.340 501.760 ;
  LAYER metal2 ;
  RECT 973.800 500.640 977.340 501.760 ;
  LAYER metal1 ;
  RECT 973.800 500.640 977.340 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 960.160 500.640 963.700 501.760 ;
  LAYER metal4 ;
  RECT 960.160 500.640 963.700 501.760 ;
  LAYER metal3 ;
  RECT 960.160 500.640 963.700 501.760 ;
  LAYER metal2 ;
  RECT 960.160 500.640 963.700 501.760 ;
  LAYER metal1 ;
  RECT 960.160 500.640 963.700 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 946.520 500.640 950.060 501.760 ;
  LAYER metal4 ;
  RECT 946.520 500.640 950.060 501.760 ;
  LAYER metal3 ;
  RECT 946.520 500.640 950.060 501.760 ;
  LAYER metal2 ;
  RECT 946.520 500.640 950.060 501.760 ;
  LAYER metal1 ;
  RECT 946.520 500.640 950.060 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 879.560 500.640 883.100 501.760 ;
  LAYER metal4 ;
  RECT 879.560 500.640 883.100 501.760 ;
  LAYER metal3 ;
  RECT 879.560 500.640 883.100 501.760 ;
  LAYER metal2 ;
  RECT 879.560 500.640 883.100 501.760 ;
  LAYER metal1 ;
  RECT 879.560 500.640 883.100 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 865.920 500.640 869.460 501.760 ;
  LAYER metal4 ;
  RECT 865.920 500.640 869.460 501.760 ;
  LAYER metal3 ;
  RECT 865.920 500.640 869.460 501.760 ;
  LAYER metal2 ;
  RECT 865.920 500.640 869.460 501.760 ;
  LAYER metal1 ;
  RECT 865.920 500.640 869.460 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 852.280 500.640 855.820 501.760 ;
  LAYER metal4 ;
  RECT 852.280 500.640 855.820 501.760 ;
  LAYER metal3 ;
  RECT 852.280 500.640 855.820 501.760 ;
  LAYER metal2 ;
  RECT 852.280 500.640 855.820 501.760 ;
  LAYER metal1 ;
  RECT 852.280 500.640 855.820 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 839.260 500.640 842.800 501.760 ;
  LAYER metal4 ;
  RECT 839.260 500.640 842.800 501.760 ;
  LAYER metal3 ;
  RECT 839.260 500.640 842.800 501.760 ;
  LAYER metal2 ;
  RECT 839.260 500.640 842.800 501.760 ;
  LAYER metal1 ;
  RECT 839.260 500.640 842.800 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 825.620 500.640 829.160 501.760 ;
  LAYER metal4 ;
  RECT 825.620 500.640 829.160 501.760 ;
  LAYER metal3 ;
  RECT 825.620 500.640 829.160 501.760 ;
  LAYER metal2 ;
  RECT 825.620 500.640 829.160 501.760 ;
  LAYER metal1 ;
  RECT 825.620 500.640 829.160 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 811.980 500.640 815.520 501.760 ;
  LAYER metal4 ;
  RECT 811.980 500.640 815.520 501.760 ;
  LAYER metal3 ;
  RECT 811.980 500.640 815.520 501.760 ;
  LAYER metal2 ;
  RECT 811.980 500.640 815.520 501.760 ;
  LAYER metal1 ;
  RECT 811.980 500.640 815.520 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 745.020 500.640 748.560 501.760 ;
  LAYER metal4 ;
  RECT 745.020 500.640 748.560 501.760 ;
  LAYER metal3 ;
  RECT 745.020 500.640 748.560 501.760 ;
  LAYER metal2 ;
  RECT 745.020 500.640 748.560 501.760 ;
  LAYER metal1 ;
  RECT 745.020 500.640 748.560 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 731.380 500.640 734.920 501.760 ;
  LAYER metal4 ;
  RECT 731.380 500.640 734.920 501.760 ;
  LAYER metal3 ;
  RECT 731.380 500.640 734.920 501.760 ;
  LAYER metal2 ;
  RECT 731.380 500.640 734.920 501.760 ;
  LAYER metal1 ;
  RECT 731.380 500.640 734.920 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 718.360 500.640 721.900 501.760 ;
  LAYER metal4 ;
  RECT 718.360 500.640 721.900 501.760 ;
  LAYER metal3 ;
  RECT 718.360 500.640 721.900 501.760 ;
  LAYER metal2 ;
  RECT 718.360 500.640 721.900 501.760 ;
  LAYER metal1 ;
  RECT 718.360 500.640 721.900 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 704.720 500.640 708.260 501.760 ;
  LAYER metal4 ;
  RECT 704.720 500.640 708.260 501.760 ;
  LAYER metal3 ;
  RECT 704.720 500.640 708.260 501.760 ;
  LAYER metal2 ;
  RECT 704.720 500.640 708.260 501.760 ;
  LAYER metal1 ;
  RECT 704.720 500.640 708.260 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 691.080 500.640 694.620 501.760 ;
  LAYER metal4 ;
  RECT 691.080 500.640 694.620 501.760 ;
  LAYER metal3 ;
  RECT 691.080 500.640 694.620 501.760 ;
  LAYER metal2 ;
  RECT 691.080 500.640 694.620 501.760 ;
  LAYER metal1 ;
  RECT 691.080 500.640 694.620 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 678.060 500.640 681.600 501.760 ;
  LAYER metal4 ;
  RECT 678.060 500.640 681.600 501.760 ;
  LAYER metal3 ;
  RECT 678.060 500.640 681.600 501.760 ;
  LAYER metal2 ;
  RECT 678.060 500.640 681.600 501.760 ;
  LAYER metal1 ;
  RECT 678.060 500.640 681.600 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 610.480 500.640 614.020 501.760 ;
  LAYER metal4 ;
  RECT 610.480 500.640 614.020 501.760 ;
  LAYER metal3 ;
  RECT 610.480 500.640 614.020 501.760 ;
  LAYER metal2 ;
  RECT 610.480 500.640 614.020 501.760 ;
  LAYER metal1 ;
  RECT 610.480 500.640 614.020 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 597.460 500.640 601.000 501.760 ;
  LAYER metal4 ;
  RECT 597.460 500.640 601.000 501.760 ;
  LAYER metal3 ;
  RECT 597.460 500.640 601.000 501.760 ;
  LAYER metal2 ;
  RECT 597.460 500.640 601.000 501.760 ;
  LAYER metal1 ;
  RECT 597.460 500.640 601.000 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 583.820 500.640 587.360 501.760 ;
  LAYER metal4 ;
  RECT 583.820 500.640 587.360 501.760 ;
  LAYER metal3 ;
  RECT 583.820 500.640 587.360 501.760 ;
  LAYER metal2 ;
  RECT 583.820 500.640 587.360 501.760 ;
  LAYER metal1 ;
  RECT 583.820 500.640 587.360 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 570.180 500.640 573.720 501.760 ;
  LAYER metal4 ;
  RECT 570.180 500.640 573.720 501.760 ;
  LAYER metal3 ;
  RECT 570.180 500.640 573.720 501.760 ;
  LAYER metal2 ;
  RECT 570.180 500.640 573.720 501.760 ;
  LAYER metal1 ;
  RECT 570.180 500.640 573.720 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 557.160 500.640 560.700 501.760 ;
  LAYER metal4 ;
  RECT 557.160 500.640 560.700 501.760 ;
  LAYER metal3 ;
  RECT 557.160 500.640 560.700 501.760 ;
  LAYER metal2 ;
  RECT 557.160 500.640 560.700 501.760 ;
  LAYER metal1 ;
  RECT 557.160 500.640 560.700 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 543.520 500.640 547.060 501.760 ;
  LAYER metal4 ;
  RECT 543.520 500.640 547.060 501.760 ;
  LAYER metal3 ;
  RECT 543.520 500.640 547.060 501.760 ;
  LAYER metal2 ;
  RECT 543.520 500.640 547.060 501.760 ;
  LAYER metal1 ;
  RECT 543.520 500.640 547.060 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 475.940 500.640 479.480 501.760 ;
  LAYER metal4 ;
  RECT 475.940 500.640 479.480 501.760 ;
  LAYER metal3 ;
  RECT 475.940 500.640 479.480 501.760 ;
  LAYER metal2 ;
  RECT 475.940 500.640 479.480 501.760 ;
  LAYER metal1 ;
  RECT 475.940 500.640 479.480 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 462.920 500.640 466.460 501.760 ;
  LAYER metal4 ;
  RECT 462.920 500.640 466.460 501.760 ;
  LAYER metal3 ;
  RECT 462.920 500.640 466.460 501.760 ;
  LAYER metal2 ;
  RECT 462.920 500.640 466.460 501.760 ;
  LAYER metal1 ;
  RECT 462.920 500.640 466.460 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 449.280 500.640 452.820 501.760 ;
  LAYER metal4 ;
  RECT 449.280 500.640 452.820 501.760 ;
  LAYER metal3 ;
  RECT 449.280 500.640 452.820 501.760 ;
  LAYER metal2 ;
  RECT 449.280 500.640 452.820 501.760 ;
  LAYER metal1 ;
  RECT 449.280 500.640 452.820 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 435.640 500.640 439.180 501.760 ;
  LAYER metal4 ;
  RECT 435.640 500.640 439.180 501.760 ;
  LAYER metal3 ;
  RECT 435.640 500.640 439.180 501.760 ;
  LAYER metal2 ;
  RECT 435.640 500.640 439.180 501.760 ;
  LAYER metal1 ;
  RECT 435.640 500.640 439.180 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 422.620 500.640 426.160 501.760 ;
  LAYER metal4 ;
  RECT 422.620 500.640 426.160 501.760 ;
  LAYER metal3 ;
  RECT 422.620 500.640 426.160 501.760 ;
  LAYER metal2 ;
  RECT 422.620 500.640 426.160 501.760 ;
  LAYER metal1 ;
  RECT 422.620 500.640 426.160 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 408.980 500.640 412.520 501.760 ;
  LAYER metal4 ;
  RECT 408.980 500.640 412.520 501.760 ;
  LAYER metal3 ;
  RECT 408.980 500.640 412.520 501.760 ;
  LAYER metal2 ;
  RECT 408.980 500.640 412.520 501.760 ;
  LAYER metal1 ;
  RECT 408.980 500.640 412.520 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 342.020 500.640 345.560 501.760 ;
  LAYER metal4 ;
  RECT 342.020 500.640 345.560 501.760 ;
  LAYER metal3 ;
  RECT 342.020 500.640 345.560 501.760 ;
  LAYER metal2 ;
  RECT 342.020 500.640 345.560 501.760 ;
  LAYER metal1 ;
  RECT 342.020 500.640 345.560 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 328.380 500.640 331.920 501.760 ;
  LAYER metal4 ;
  RECT 328.380 500.640 331.920 501.760 ;
  LAYER metal3 ;
  RECT 328.380 500.640 331.920 501.760 ;
  LAYER metal2 ;
  RECT 328.380 500.640 331.920 501.760 ;
  LAYER metal1 ;
  RECT 328.380 500.640 331.920 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 314.740 500.640 318.280 501.760 ;
  LAYER metal4 ;
  RECT 314.740 500.640 318.280 501.760 ;
  LAYER metal3 ;
  RECT 314.740 500.640 318.280 501.760 ;
  LAYER metal2 ;
  RECT 314.740 500.640 318.280 501.760 ;
  LAYER metal1 ;
  RECT 314.740 500.640 318.280 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 301.720 500.640 305.260 501.760 ;
  LAYER metal4 ;
  RECT 301.720 500.640 305.260 501.760 ;
  LAYER metal3 ;
  RECT 301.720 500.640 305.260 501.760 ;
  LAYER metal2 ;
  RECT 301.720 500.640 305.260 501.760 ;
  LAYER metal1 ;
  RECT 301.720 500.640 305.260 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 288.080 500.640 291.620 501.760 ;
  LAYER metal4 ;
  RECT 288.080 500.640 291.620 501.760 ;
  LAYER metal3 ;
  RECT 288.080 500.640 291.620 501.760 ;
  LAYER metal2 ;
  RECT 288.080 500.640 291.620 501.760 ;
  LAYER metal1 ;
  RECT 288.080 500.640 291.620 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 274.440 500.640 277.980 501.760 ;
  LAYER metal4 ;
  RECT 274.440 500.640 277.980 501.760 ;
  LAYER metal3 ;
  RECT 274.440 500.640 277.980 501.760 ;
  LAYER metal2 ;
  RECT 274.440 500.640 277.980 501.760 ;
  LAYER metal1 ;
  RECT 274.440 500.640 277.980 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 207.480 500.640 211.020 501.760 ;
  LAYER metal4 ;
  RECT 207.480 500.640 211.020 501.760 ;
  LAYER metal3 ;
  RECT 207.480 500.640 211.020 501.760 ;
  LAYER metal2 ;
  RECT 207.480 500.640 211.020 501.760 ;
  LAYER metal1 ;
  RECT 207.480 500.640 211.020 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 193.840 500.640 197.380 501.760 ;
  LAYER metal4 ;
  RECT 193.840 500.640 197.380 501.760 ;
  LAYER metal3 ;
  RECT 193.840 500.640 197.380 501.760 ;
  LAYER metal2 ;
  RECT 193.840 500.640 197.380 501.760 ;
  LAYER metal1 ;
  RECT 193.840 500.640 197.380 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 180.820 500.640 184.360 501.760 ;
  LAYER metal4 ;
  RECT 180.820 500.640 184.360 501.760 ;
  LAYER metal3 ;
  RECT 180.820 500.640 184.360 501.760 ;
  LAYER metal2 ;
  RECT 180.820 500.640 184.360 501.760 ;
  LAYER metal1 ;
  RECT 180.820 500.640 184.360 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 167.180 500.640 170.720 501.760 ;
  LAYER metal4 ;
  RECT 167.180 500.640 170.720 501.760 ;
  LAYER metal3 ;
  RECT 167.180 500.640 170.720 501.760 ;
  LAYER metal2 ;
  RECT 167.180 500.640 170.720 501.760 ;
  LAYER metal1 ;
  RECT 167.180 500.640 170.720 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 153.540 500.640 157.080 501.760 ;
  LAYER metal4 ;
  RECT 153.540 500.640 157.080 501.760 ;
  LAYER metal3 ;
  RECT 153.540 500.640 157.080 501.760 ;
  LAYER metal2 ;
  RECT 153.540 500.640 157.080 501.760 ;
  LAYER metal1 ;
  RECT 153.540 500.640 157.080 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 140.520 500.640 144.060 501.760 ;
  LAYER metal4 ;
  RECT 140.520 500.640 144.060 501.760 ;
  LAYER metal3 ;
  RECT 140.520 500.640 144.060 501.760 ;
  LAYER metal2 ;
  RECT 140.520 500.640 144.060 501.760 ;
  LAYER metal1 ;
  RECT 140.520 500.640 144.060 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 72.940 500.640 76.480 501.760 ;
  LAYER metal4 ;
  RECT 72.940 500.640 76.480 501.760 ;
  LAYER metal3 ;
  RECT 72.940 500.640 76.480 501.760 ;
  LAYER metal2 ;
  RECT 72.940 500.640 76.480 501.760 ;
  LAYER metal1 ;
  RECT 72.940 500.640 76.480 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 59.300 500.640 62.840 501.760 ;
  LAYER metal4 ;
  RECT 59.300 500.640 62.840 501.760 ;
  LAYER metal3 ;
  RECT 59.300 500.640 62.840 501.760 ;
  LAYER metal2 ;
  RECT 59.300 500.640 62.840 501.760 ;
  LAYER metal1 ;
  RECT 59.300 500.640 62.840 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 46.280 500.640 49.820 501.760 ;
  LAYER metal4 ;
  RECT 46.280 500.640 49.820 501.760 ;
  LAYER metal3 ;
  RECT 46.280 500.640 49.820 501.760 ;
  LAYER metal2 ;
  RECT 46.280 500.640 49.820 501.760 ;
  LAYER metal1 ;
  RECT 46.280 500.640 49.820 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 32.640 500.640 36.180 501.760 ;
  LAYER metal4 ;
  RECT 32.640 500.640 36.180 501.760 ;
  LAYER metal3 ;
  RECT 32.640 500.640 36.180 501.760 ;
  LAYER metal2 ;
  RECT 32.640 500.640 36.180 501.760 ;
  LAYER metal1 ;
  RECT 32.640 500.640 36.180 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 19.000 500.640 22.540 501.760 ;
  LAYER metal4 ;
  RECT 19.000 500.640 22.540 501.760 ;
  LAYER metal3 ;
  RECT 19.000 500.640 22.540 501.760 ;
  LAYER metal2 ;
  RECT 19.000 500.640 22.540 501.760 ;
  LAYER metal1 ;
  RECT 19.000 500.640 22.540 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 7.220 500.640 10.760 501.760 ;
  LAYER metal4 ;
  RECT 7.220 500.640 10.760 501.760 ;
  LAYER metal3 ;
  RECT 7.220 500.640 10.760 501.760 ;
  LAYER metal2 ;
  RECT 7.220 500.640 10.760 501.760 ;
  LAYER metal1 ;
  RECT 7.220 500.640 10.760 501.760 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3584.000 0.000 3587.540 1.120 ;
  LAYER metal4 ;
  RECT 3584.000 0.000 3587.540 1.120 ;
  LAYER metal3 ;
  RECT 3584.000 0.000 3587.540 1.120 ;
  LAYER metal2 ;
  RECT 3584.000 0.000 3587.540 1.120 ;
  LAYER metal1 ;
  RECT 3584.000 0.000 3587.540 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3575.320 0.000 3578.860 1.120 ;
  LAYER metal4 ;
  RECT 3575.320 0.000 3578.860 1.120 ;
  LAYER metal3 ;
  RECT 3575.320 0.000 3578.860 1.120 ;
  LAYER metal2 ;
  RECT 3575.320 0.000 3578.860 1.120 ;
  LAYER metal1 ;
  RECT 3575.320 0.000 3578.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3561.680 0.000 3565.220 1.120 ;
  LAYER metal4 ;
  RECT 3561.680 0.000 3565.220 1.120 ;
  LAYER metal3 ;
  RECT 3561.680 0.000 3565.220 1.120 ;
  LAYER metal2 ;
  RECT 3561.680 0.000 3565.220 1.120 ;
  LAYER metal1 ;
  RECT 3561.680 0.000 3565.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3548.660 0.000 3552.200 1.120 ;
  LAYER metal4 ;
  RECT 3548.660 0.000 3552.200 1.120 ;
  LAYER metal3 ;
  RECT 3548.660 0.000 3552.200 1.120 ;
  LAYER metal2 ;
  RECT 3548.660 0.000 3552.200 1.120 ;
  LAYER metal1 ;
  RECT 3548.660 0.000 3552.200 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3535.020 0.000 3538.560 1.120 ;
  LAYER metal4 ;
  RECT 3535.020 0.000 3538.560 1.120 ;
  LAYER metal3 ;
  RECT 3535.020 0.000 3538.560 1.120 ;
  LAYER metal2 ;
  RECT 3535.020 0.000 3538.560 1.120 ;
  LAYER metal1 ;
  RECT 3535.020 0.000 3538.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3521.380 0.000 3524.920 1.120 ;
  LAYER metal4 ;
  RECT 3521.380 0.000 3524.920 1.120 ;
  LAYER metal3 ;
  RECT 3521.380 0.000 3524.920 1.120 ;
  LAYER metal2 ;
  RECT 3521.380 0.000 3524.920 1.120 ;
  LAYER metal1 ;
  RECT 3521.380 0.000 3524.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3454.420 0.000 3457.960 1.120 ;
  LAYER metal4 ;
  RECT 3454.420 0.000 3457.960 1.120 ;
  LAYER metal3 ;
  RECT 3454.420 0.000 3457.960 1.120 ;
  LAYER metal2 ;
  RECT 3454.420 0.000 3457.960 1.120 ;
  LAYER metal1 ;
  RECT 3454.420 0.000 3457.960 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3440.780 0.000 3444.320 1.120 ;
  LAYER metal4 ;
  RECT 3440.780 0.000 3444.320 1.120 ;
  LAYER metal3 ;
  RECT 3440.780 0.000 3444.320 1.120 ;
  LAYER metal2 ;
  RECT 3440.780 0.000 3444.320 1.120 ;
  LAYER metal1 ;
  RECT 3440.780 0.000 3444.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3427.760 0.000 3431.300 1.120 ;
  LAYER metal4 ;
  RECT 3427.760 0.000 3431.300 1.120 ;
  LAYER metal3 ;
  RECT 3427.760 0.000 3431.300 1.120 ;
  LAYER metal2 ;
  RECT 3427.760 0.000 3431.300 1.120 ;
  LAYER metal1 ;
  RECT 3427.760 0.000 3431.300 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3414.120 0.000 3417.660 1.120 ;
  LAYER metal4 ;
  RECT 3414.120 0.000 3417.660 1.120 ;
  LAYER metal3 ;
  RECT 3414.120 0.000 3417.660 1.120 ;
  LAYER metal2 ;
  RECT 3414.120 0.000 3417.660 1.120 ;
  LAYER metal1 ;
  RECT 3414.120 0.000 3417.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3400.480 0.000 3404.020 1.120 ;
  LAYER metal4 ;
  RECT 3400.480 0.000 3404.020 1.120 ;
  LAYER metal3 ;
  RECT 3400.480 0.000 3404.020 1.120 ;
  LAYER metal2 ;
  RECT 3400.480 0.000 3404.020 1.120 ;
  LAYER metal1 ;
  RECT 3400.480 0.000 3404.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3387.460 0.000 3391.000 1.120 ;
  LAYER metal4 ;
  RECT 3387.460 0.000 3391.000 1.120 ;
  LAYER metal3 ;
  RECT 3387.460 0.000 3391.000 1.120 ;
  LAYER metal2 ;
  RECT 3387.460 0.000 3391.000 1.120 ;
  LAYER metal1 ;
  RECT 3387.460 0.000 3391.000 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3319.880 0.000 3323.420 1.120 ;
  LAYER metal4 ;
  RECT 3319.880 0.000 3323.420 1.120 ;
  LAYER metal3 ;
  RECT 3319.880 0.000 3323.420 1.120 ;
  LAYER metal2 ;
  RECT 3319.880 0.000 3323.420 1.120 ;
  LAYER metal1 ;
  RECT 3319.880 0.000 3323.420 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3306.860 0.000 3310.400 1.120 ;
  LAYER metal4 ;
  RECT 3306.860 0.000 3310.400 1.120 ;
  LAYER metal3 ;
  RECT 3306.860 0.000 3310.400 1.120 ;
  LAYER metal2 ;
  RECT 3306.860 0.000 3310.400 1.120 ;
  LAYER metal1 ;
  RECT 3306.860 0.000 3310.400 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3293.220 0.000 3296.760 1.120 ;
  LAYER metal4 ;
  RECT 3293.220 0.000 3296.760 1.120 ;
  LAYER metal3 ;
  RECT 3293.220 0.000 3296.760 1.120 ;
  LAYER metal2 ;
  RECT 3293.220 0.000 3296.760 1.120 ;
  LAYER metal1 ;
  RECT 3293.220 0.000 3296.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3279.580 0.000 3283.120 1.120 ;
  LAYER metal4 ;
  RECT 3279.580 0.000 3283.120 1.120 ;
  LAYER metal3 ;
  RECT 3279.580 0.000 3283.120 1.120 ;
  LAYER metal2 ;
  RECT 3279.580 0.000 3283.120 1.120 ;
  LAYER metal1 ;
  RECT 3279.580 0.000 3283.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3266.560 0.000 3270.100 1.120 ;
  LAYER metal4 ;
  RECT 3266.560 0.000 3270.100 1.120 ;
  LAYER metal3 ;
  RECT 3266.560 0.000 3270.100 1.120 ;
  LAYER metal2 ;
  RECT 3266.560 0.000 3270.100 1.120 ;
  LAYER metal1 ;
  RECT 3266.560 0.000 3270.100 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3252.920 0.000 3256.460 1.120 ;
  LAYER metal4 ;
  RECT 3252.920 0.000 3256.460 1.120 ;
  LAYER metal3 ;
  RECT 3252.920 0.000 3256.460 1.120 ;
  LAYER metal2 ;
  RECT 3252.920 0.000 3256.460 1.120 ;
  LAYER metal1 ;
  RECT 3252.920 0.000 3256.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3185.960 0.000 3189.500 1.120 ;
  LAYER metal4 ;
  RECT 3185.960 0.000 3189.500 1.120 ;
  LAYER metal3 ;
  RECT 3185.960 0.000 3189.500 1.120 ;
  LAYER metal2 ;
  RECT 3185.960 0.000 3189.500 1.120 ;
  LAYER metal1 ;
  RECT 3185.960 0.000 3189.500 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3172.320 0.000 3175.860 1.120 ;
  LAYER metal4 ;
  RECT 3172.320 0.000 3175.860 1.120 ;
  LAYER metal3 ;
  RECT 3172.320 0.000 3175.860 1.120 ;
  LAYER metal2 ;
  RECT 3172.320 0.000 3175.860 1.120 ;
  LAYER metal1 ;
  RECT 3172.320 0.000 3175.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3158.680 0.000 3162.220 1.120 ;
  LAYER metal4 ;
  RECT 3158.680 0.000 3162.220 1.120 ;
  LAYER metal3 ;
  RECT 3158.680 0.000 3162.220 1.120 ;
  LAYER metal2 ;
  RECT 3158.680 0.000 3162.220 1.120 ;
  LAYER metal1 ;
  RECT 3158.680 0.000 3162.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3145.040 0.000 3148.580 1.120 ;
  LAYER metal4 ;
  RECT 3145.040 0.000 3148.580 1.120 ;
  LAYER metal3 ;
  RECT 3145.040 0.000 3148.580 1.120 ;
  LAYER metal2 ;
  RECT 3145.040 0.000 3148.580 1.120 ;
  LAYER metal1 ;
  RECT 3145.040 0.000 3148.580 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3132.020 0.000 3135.560 1.120 ;
  LAYER metal4 ;
  RECT 3132.020 0.000 3135.560 1.120 ;
  LAYER metal3 ;
  RECT 3132.020 0.000 3135.560 1.120 ;
  LAYER metal2 ;
  RECT 3132.020 0.000 3135.560 1.120 ;
  LAYER metal1 ;
  RECT 3132.020 0.000 3135.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3118.380 0.000 3121.920 1.120 ;
  LAYER metal4 ;
  RECT 3118.380 0.000 3121.920 1.120 ;
  LAYER metal3 ;
  RECT 3118.380 0.000 3121.920 1.120 ;
  LAYER metal2 ;
  RECT 3118.380 0.000 3121.920 1.120 ;
  LAYER metal1 ;
  RECT 3118.380 0.000 3121.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3051.420 0.000 3054.960 1.120 ;
  LAYER metal4 ;
  RECT 3051.420 0.000 3054.960 1.120 ;
  LAYER metal3 ;
  RECT 3051.420 0.000 3054.960 1.120 ;
  LAYER metal2 ;
  RECT 3051.420 0.000 3054.960 1.120 ;
  LAYER metal1 ;
  RECT 3051.420 0.000 3054.960 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3037.780 0.000 3041.320 1.120 ;
  LAYER metal4 ;
  RECT 3037.780 0.000 3041.320 1.120 ;
  LAYER metal3 ;
  RECT 3037.780 0.000 3041.320 1.120 ;
  LAYER metal2 ;
  RECT 3037.780 0.000 3041.320 1.120 ;
  LAYER metal1 ;
  RECT 3037.780 0.000 3041.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3024.140 0.000 3027.680 1.120 ;
  LAYER metal4 ;
  RECT 3024.140 0.000 3027.680 1.120 ;
  LAYER metal3 ;
  RECT 3024.140 0.000 3027.680 1.120 ;
  LAYER metal2 ;
  RECT 3024.140 0.000 3027.680 1.120 ;
  LAYER metal1 ;
  RECT 3024.140 0.000 3027.680 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3011.120 0.000 3014.660 1.120 ;
  LAYER metal4 ;
  RECT 3011.120 0.000 3014.660 1.120 ;
  LAYER metal3 ;
  RECT 3011.120 0.000 3014.660 1.120 ;
  LAYER metal2 ;
  RECT 3011.120 0.000 3014.660 1.120 ;
  LAYER metal1 ;
  RECT 3011.120 0.000 3014.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2997.480 0.000 3001.020 1.120 ;
  LAYER metal4 ;
  RECT 2997.480 0.000 3001.020 1.120 ;
  LAYER metal3 ;
  RECT 2997.480 0.000 3001.020 1.120 ;
  LAYER metal2 ;
  RECT 2997.480 0.000 3001.020 1.120 ;
  LAYER metal1 ;
  RECT 2997.480 0.000 3001.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2983.840 0.000 2987.380 1.120 ;
  LAYER metal4 ;
  RECT 2983.840 0.000 2987.380 1.120 ;
  LAYER metal3 ;
  RECT 2983.840 0.000 2987.380 1.120 ;
  LAYER metal2 ;
  RECT 2983.840 0.000 2987.380 1.120 ;
  LAYER metal1 ;
  RECT 2983.840 0.000 2987.380 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2916.880 0.000 2920.420 1.120 ;
  LAYER metal4 ;
  RECT 2916.880 0.000 2920.420 1.120 ;
  LAYER metal3 ;
  RECT 2916.880 0.000 2920.420 1.120 ;
  LAYER metal2 ;
  RECT 2916.880 0.000 2920.420 1.120 ;
  LAYER metal1 ;
  RECT 2916.880 0.000 2920.420 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2903.240 0.000 2906.780 1.120 ;
  LAYER metal4 ;
  RECT 2903.240 0.000 2906.780 1.120 ;
  LAYER metal3 ;
  RECT 2903.240 0.000 2906.780 1.120 ;
  LAYER metal2 ;
  RECT 2903.240 0.000 2906.780 1.120 ;
  LAYER metal1 ;
  RECT 2903.240 0.000 2906.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2890.220 0.000 2893.760 1.120 ;
  LAYER metal4 ;
  RECT 2890.220 0.000 2893.760 1.120 ;
  LAYER metal3 ;
  RECT 2890.220 0.000 2893.760 1.120 ;
  LAYER metal2 ;
  RECT 2890.220 0.000 2893.760 1.120 ;
  LAYER metal1 ;
  RECT 2890.220 0.000 2893.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2876.580 0.000 2880.120 1.120 ;
  LAYER metal4 ;
  RECT 2876.580 0.000 2880.120 1.120 ;
  LAYER metal3 ;
  RECT 2876.580 0.000 2880.120 1.120 ;
  LAYER metal2 ;
  RECT 2876.580 0.000 2880.120 1.120 ;
  LAYER metal1 ;
  RECT 2876.580 0.000 2880.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2862.940 0.000 2866.480 1.120 ;
  LAYER metal4 ;
  RECT 2862.940 0.000 2866.480 1.120 ;
  LAYER metal3 ;
  RECT 2862.940 0.000 2866.480 1.120 ;
  LAYER metal2 ;
  RECT 2862.940 0.000 2866.480 1.120 ;
  LAYER metal1 ;
  RECT 2862.940 0.000 2866.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2849.920 0.000 2853.460 1.120 ;
  LAYER metal4 ;
  RECT 2849.920 0.000 2853.460 1.120 ;
  LAYER metal3 ;
  RECT 2849.920 0.000 2853.460 1.120 ;
  LAYER metal2 ;
  RECT 2849.920 0.000 2853.460 1.120 ;
  LAYER metal1 ;
  RECT 2849.920 0.000 2853.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2782.340 0.000 2785.880 1.120 ;
  LAYER metal4 ;
  RECT 2782.340 0.000 2785.880 1.120 ;
  LAYER metal3 ;
  RECT 2782.340 0.000 2785.880 1.120 ;
  LAYER metal2 ;
  RECT 2782.340 0.000 2785.880 1.120 ;
  LAYER metal1 ;
  RECT 2782.340 0.000 2785.880 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2769.320 0.000 2772.860 1.120 ;
  LAYER metal4 ;
  RECT 2769.320 0.000 2772.860 1.120 ;
  LAYER metal3 ;
  RECT 2769.320 0.000 2772.860 1.120 ;
  LAYER metal2 ;
  RECT 2769.320 0.000 2772.860 1.120 ;
  LAYER metal1 ;
  RECT 2769.320 0.000 2772.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2755.680 0.000 2759.220 1.120 ;
  LAYER metal4 ;
  RECT 2755.680 0.000 2759.220 1.120 ;
  LAYER metal3 ;
  RECT 2755.680 0.000 2759.220 1.120 ;
  LAYER metal2 ;
  RECT 2755.680 0.000 2759.220 1.120 ;
  LAYER metal1 ;
  RECT 2755.680 0.000 2759.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2742.040 0.000 2745.580 1.120 ;
  LAYER metal4 ;
  RECT 2742.040 0.000 2745.580 1.120 ;
  LAYER metal3 ;
  RECT 2742.040 0.000 2745.580 1.120 ;
  LAYER metal2 ;
  RECT 2742.040 0.000 2745.580 1.120 ;
  LAYER metal1 ;
  RECT 2742.040 0.000 2745.580 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2728.400 0.000 2731.940 1.120 ;
  LAYER metal4 ;
  RECT 2728.400 0.000 2731.940 1.120 ;
  LAYER metal3 ;
  RECT 2728.400 0.000 2731.940 1.120 ;
  LAYER metal2 ;
  RECT 2728.400 0.000 2731.940 1.120 ;
  LAYER metal1 ;
  RECT 2728.400 0.000 2731.940 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2715.380 0.000 2718.920 1.120 ;
  LAYER metal4 ;
  RECT 2715.380 0.000 2718.920 1.120 ;
  LAYER metal3 ;
  RECT 2715.380 0.000 2718.920 1.120 ;
  LAYER metal2 ;
  RECT 2715.380 0.000 2718.920 1.120 ;
  LAYER metal1 ;
  RECT 2715.380 0.000 2718.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2647.800 0.000 2651.340 1.120 ;
  LAYER metal4 ;
  RECT 2647.800 0.000 2651.340 1.120 ;
  LAYER metal3 ;
  RECT 2647.800 0.000 2651.340 1.120 ;
  LAYER metal2 ;
  RECT 2647.800 0.000 2651.340 1.120 ;
  LAYER metal1 ;
  RECT 2647.800 0.000 2651.340 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2634.780 0.000 2638.320 1.120 ;
  LAYER metal4 ;
  RECT 2634.780 0.000 2638.320 1.120 ;
  LAYER metal3 ;
  RECT 2634.780 0.000 2638.320 1.120 ;
  LAYER metal2 ;
  RECT 2634.780 0.000 2638.320 1.120 ;
  LAYER metal1 ;
  RECT 2634.780 0.000 2638.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2621.140 0.000 2624.680 1.120 ;
  LAYER metal4 ;
  RECT 2621.140 0.000 2624.680 1.120 ;
  LAYER metal3 ;
  RECT 2621.140 0.000 2624.680 1.120 ;
  LAYER metal2 ;
  RECT 2621.140 0.000 2624.680 1.120 ;
  LAYER metal1 ;
  RECT 2621.140 0.000 2624.680 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2607.500 0.000 2611.040 1.120 ;
  LAYER metal4 ;
  RECT 2607.500 0.000 2611.040 1.120 ;
  LAYER metal3 ;
  RECT 2607.500 0.000 2611.040 1.120 ;
  LAYER metal2 ;
  RECT 2607.500 0.000 2611.040 1.120 ;
  LAYER metal1 ;
  RECT 2607.500 0.000 2611.040 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2594.480 0.000 2598.020 1.120 ;
  LAYER metal4 ;
  RECT 2594.480 0.000 2598.020 1.120 ;
  LAYER metal3 ;
  RECT 2594.480 0.000 2598.020 1.120 ;
  LAYER metal2 ;
  RECT 2594.480 0.000 2598.020 1.120 ;
  LAYER metal1 ;
  RECT 2594.480 0.000 2598.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2580.840 0.000 2584.380 1.120 ;
  LAYER metal4 ;
  RECT 2580.840 0.000 2584.380 1.120 ;
  LAYER metal3 ;
  RECT 2580.840 0.000 2584.380 1.120 ;
  LAYER metal2 ;
  RECT 2580.840 0.000 2584.380 1.120 ;
  LAYER metal1 ;
  RECT 2580.840 0.000 2584.380 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2513.880 0.000 2517.420 1.120 ;
  LAYER metal4 ;
  RECT 2513.880 0.000 2517.420 1.120 ;
  LAYER metal3 ;
  RECT 2513.880 0.000 2517.420 1.120 ;
  LAYER metal2 ;
  RECT 2513.880 0.000 2517.420 1.120 ;
  LAYER metal1 ;
  RECT 2513.880 0.000 2517.420 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2500.240 0.000 2503.780 1.120 ;
  LAYER metal4 ;
  RECT 2500.240 0.000 2503.780 1.120 ;
  LAYER metal3 ;
  RECT 2500.240 0.000 2503.780 1.120 ;
  LAYER metal2 ;
  RECT 2500.240 0.000 2503.780 1.120 ;
  LAYER metal1 ;
  RECT 2500.240 0.000 2503.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2486.600 0.000 2490.140 1.120 ;
  LAYER metal4 ;
  RECT 2486.600 0.000 2490.140 1.120 ;
  LAYER metal3 ;
  RECT 2486.600 0.000 2490.140 1.120 ;
  LAYER metal2 ;
  RECT 2486.600 0.000 2490.140 1.120 ;
  LAYER metal1 ;
  RECT 2486.600 0.000 2490.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2473.580 0.000 2477.120 1.120 ;
  LAYER metal4 ;
  RECT 2473.580 0.000 2477.120 1.120 ;
  LAYER metal3 ;
  RECT 2473.580 0.000 2477.120 1.120 ;
  LAYER metal2 ;
  RECT 2473.580 0.000 2477.120 1.120 ;
  LAYER metal1 ;
  RECT 2473.580 0.000 2477.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2459.940 0.000 2463.480 1.120 ;
  LAYER metal4 ;
  RECT 2459.940 0.000 2463.480 1.120 ;
  LAYER metal3 ;
  RECT 2459.940 0.000 2463.480 1.120 ;
  LAYER metal2 ;
  RECT 2459.940 0.000 2463.480 1.120 ;
  LAYER metal1 ;
  RECT 2459.940 0.000 2463.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2446.300 0.000 2449.840 1.120 ;
  LAYER metal4 ;
  RECT 2446.300 0.000 2449.840 1.120 ;
  LAYER metal3 ;
  RECT 2446.300 0.000 2449.840 1.120 ;
  LAYER metal2 ;
  RECT 2446.300 0.000 2449.840 1.120 ;
  LAYER metal1 ;
  RECT 2446.300 0.000 2449.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2379.340 0.000 2382.880 1.120 ;
  LAYER metal4 ;
  RECT 2379.340 0.000 2382.880 1.120 ;
  LAYER metal3 ;
  RECT 2379.340 0.000 2382.880 1.120 ;
  LAYER metal2 ;
  RECT 2379.340 0.000 2382.880 1.120 ;
  LAYER metal1 ;
  RECT 2379.340 0.000 2382.880 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2365.700 0.000 2369.240 1.120 ;
  LAYER metal4 ;
  RECT 2365.700 0.000 2369.240 1.120 ;
  LAYER metal3 ;
  RECT 2365.700 0.000 2369.240 1.120 ;
  LAYER metal2 ;
  RECT 2365.700 0.000 2369.240 1.120 ;
  LAYER metal1 ;
  RECT 2365.700 0.000 2369.240 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2352.680 0.000 2356.220 1.120 ;
  LAYER metal4 ;
  RECT 2352.680 0.000 2356.220 1.120 ;
  LAYER metal3 ;
  RECT 2352.680 0.000 2356.220 1.120 ;
  LAYER metal2 ;
  RECT 2352.680 0.000 2356.220 1.120 ;
  LAYER metal1 ;
  RECT 2352.680 0.000 2356.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2339.040 0.000 2342.580 1.120 ;
  LAYER metal4 ;
  RECT 2339.040 0.000 2342.580 1.120 ;
  LAYER metal3 ;
  RECT 2339.040 0.000 2342.580 1.120 ;
  LAYER metal2 ;
  RECT 2339.040 0.000 2342.580 1.120 ;
  LAYER metal1 ;
  RECT 2339.040 0.000 2342.580 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2325.400 0.000 2328.940 1.120 ;
  LAYER metal4 ;
  RECT 2325.400 0.000 2328.940 1.120 ;
  LAYER metal3 ;
  RECT 2325.400 0.000 2328.940 1.120 ;
  LAYER metal2 ;
  RECT 2325.400 0.000 2328.940 1.120 ;
  LAYER metal1 ;
  RECT 2325.400 0.000 2328.940 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2311.760 0.000 2315.300 1.120 ;
  LAYER metal4 ;
  RECT 2311.760 0.000 2315.300 1.120 ;
  LAYER metal3 ;
  RECT 2311.760 0.000 2315.300 1.120 ;
  LAYER metal2 ;
  RECT 2311.760 0.000 2315.300 1.120 ;
  LAYER metal1 ;
  RECT 2311.760 0.000 2315.300 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2244.800 0.000 2248.340 1.120 ;
  LAYER metal4 ;
  RECT 2244.800 0.000 2248.340 1.120 ;
  LAYER metal3 ;
  RECT 2244.800 0.000 2248.340 1.120 ;
  LAYER metal2 ;
  RECT 2244.800 0.000 2248.340 1.120 ;
  LAYER metal1 ;
  RECT 2244.800 0.000 2248.340 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2231.160 0.000 2234.700 1.120 ;
  LAYER metal4 ;
  RECT 2231.160 0.000 2234.700 1.120 ;
  LAYER metal3 ;
  RECT 2231.160 0.000 2234.700 1.120 ;
  LAYER metal2 ;
  RECT 2231.160 0.000 2234.700 1.120 ;
  LAYER metal1 ;
  RECT 2231.160 0.000 2234.700 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2218.140 0.000 2221.680 1.120 ;
  LAYER metal4 ;
  RECT 2218.140 0.000 2221.680 1.120 ;
  LAYER metal3 ;
  RECT 2218.140 0.000 2221.680 1.120 ;
  LAYER metal2 ;
  RECT 2218.140 0.000 2221.680 1.120 ;
  LAYER metal1 ;
  RECT 2218.140 0.000 2221.680 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2204.500 0.000 2208.040 1.120 ;
  LAYER metal4 ;
  RECT 2204.500 0.000 2208.040 1.120 ;
  LAYER metal3 ;
  RECT 2204.500 0.000 2208.040 1.120 ;
  LAYER metal2 ;
  RECT 2204.500 0.000 2208.040 1.120 ;
  LAYER metal1 ;
  RECT 2204.500 0.000 2208.040 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2190.860 0.000 2194.400 1.120 ;
  LAYER metal4 ;
  RECT 2190.860 0.000 2194.400 1.120 ;
  LAYER metal3 ;
  RECT 2190.860 0.000 2194.400 1.120 ;
  LAYER metal2 ;
  RECT 2190.860 0.000 2194.400 1.120 ;
  LAYER metal1 ;
  RECT 2190.860 0.000 2194.400 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2177.840 0.000 2181.380 1.120 ;
  LAYER metal4 ;
  RECT 2177.840 0.000 2181.380 1.120 ;
  LAYER metal3 ;
  RECT 2177.840 0.000 2181.380 1.120 ;
  LAYER metal2 ;
  RECT 2177.840 0.000 2181.380 1.120 ;
  LAYER metal1 ;
  RECT 2177.840 0.000 2181.380 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2110.260 0.000 2113.800 1.120 ;
  LAYER metal4 ;
  RECT 2110.260 0.000 2113.800 1.120 ;
  LAYER metal3 ;
  RECT 2110.260 0.000 2113.800 1.120 ;
  LAYER metal2 ;
  RECT 2110.260 0.000 2113.800 1.120 ;
  LAYER metal1 ;
  RECT 2110.260 0.000 2113.800 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2097.240 0.000 2100.780 1.120 ;
  LAYER metal4 ;
  RECT 2097.240 0.000 2100.780 1.120 ;
  LAYER metal3 ;
  RECT 2097.240 0.000 2100.780 1.120 ;
  LAYER metal2 ;
  RECT 2097.240 0.000 2100.780 1.120 ;
  LAYER metal1 ;
  RECT 2097.240 0.000 2100.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2083.600 0.000 2087.140 1.120 ;
  LAYER metal4 ;
  RECT 2083.600 0.000 2087.140 1.120 ;
  LAYER metal3 ;
  RECT 2083.600 0.000 2087.140 1.120 ;
  LAYER metal2 ;
  RECT 2083.600 0.000 2087.140 1.120 ;
  LAYER metal1 ;
  RECT 2083.600 0.000 2087.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2069.960 0.000 2073.500 1.120 ;
  LAYER metal4 ;
  RECT 2069.960 0.000 2073.500 1.120 ;
  LAYER metal3 ;
  RECT 2069.960 0.000 2073.500 1.120 ;
  LAYER metal2 ;
  RECT 2069.960 0.000 2073.500 1.120 ;
  LAYER metal1 ;
  RECT 2069.960 0.000 2073.500 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2056.940 0.000 2060.480 1.120 ;
  LAYER metal4 ;
  RECT 2056.940 0.000 2060.480 1.120 ;
  LAYER metal3 ;
  RECT 2056.940 0.000 2060.480 1.120 ;
  LAYER metal2 ;
  RECT 2056.940 0.000 2060.480 1.120 ;
  LAYER metal1 ;
  RECT 2056.940 0.000 2060.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2043.300 0.000 2046.840 1.120 ;
  LAYER metal4 ;
  RECT 2043.300 0.000 2046.840 1.120 ;
  LAYER metal3 ;
  RECT 2043.300 0.000 2046.840 1.120 ;
  LAYER metal2 ;
  RECT 2043.300 0.000 2046.840 1.120 ;
  LAYER metal1 ;
  RECT 2043.300 0.000 2046.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1976.340 0.000 1979.880 1.120 ;
  LAYER metal4 ;
  RECT 1976.340 0.000 1979.880 1.120 ;
  LAYER metal3 ;
  RECT 1976.340 0.000 1979.880 1.120 ;
  LAYER metal2 ;
  RECT 1976.340 0.000 1979.880 1.120 ;
  LAYER metal1 ;
  RECT 1976.340 0.000 1979.880 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1962.700 0.000 1966.240 1.120 ;
  LAYER metal4 ;
  RECT 1962.700 0.000 1966.240 1.120 ;
  LAYER metal3 ;
  RECT 1962.700 0.000 1966.240 1.120 ;
  LAYER metal2 ;
  RECT 1962.700 0.000 1966.240 1.120 ;
  LAYER metal1 ;
  RECT 1962.700 0.000 1966.240 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1949.060 0.000 1952.600 1.120 ;
  LAYER metal4 ;
  RECT 1949.060 0.000 1952.600 1.120 ;
  LAYER metal3 ;
  RECT 1949.060 0.000 1952.600 1.120 ;
  LAYER metal2 ;
  RECT 1949.060 0.000 1952.600 1.120 ;
  LAYER metal1 ;
  RECT 1949.060 0.000 1952.600 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1936.040 0.000 1939.580 1.120 ;
  LAYER metal4 ;
  RECT 1936.040 0.000 1939.580 1.120 ;
  LAYER metal3 ;
  RECT 1936.040 0.000 1939.580 1.120 ;
  LAYER metal2 ;
  RECT 1936.040 0.000 1939.580 1.120 ;
  LAYER metal1 ;
  RECT 1936.040 0.000 1939.580 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1922.400 0.000 1925.940 1.120 ;
  LAYER metal4 ;
  RECT 1922.400 0.000 1925.940 1.120 ;
  LAYER metal3 ;
  RECT 1922.400 0.000 1925.940 1.120 ;
  LAYER metal2 ;
  RECT 1922.400 0.000 1925.940 1.120 ;
  LAYER metal1 ;
  RECT 1922.400 0.000 1925.940 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1908.760 0.000 1912.300 1.120 ;
  LAYER metal4 ;
  RECT 1908.760 0.000 1912.300 1.120 ;
  LAYER metal3 ;
  RECT 1908.760 0.000 1912.300 1.120 ;
  LAYER metal2 ;
  RECT 1908.760 0.000 1912.300 1.120 ;
  LAYER metal1 ;
  RECT 1908.760 0.000 1912.300 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1846.140 0.000 1849.680 1.120 ;
  LAYER metal4 ;
  RECT 1846.140 0.000 1849.680 1.120 ;
  LAYER metal3 ;
  RECT 1846.140 0.000 1849.680 1.120 ;
  LAYER metal2 ;
  RECT 1846.140 0.000 1849.680 1.120 ;
  LAYER metal1 ;
  RECT 1846.140 0.000 1849.680 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1833.120 0.000 1836.660 1.120 ;
  LAYER metal4 ;
  RECT 1833.120 0.000 1836.660 1.120 ;
  LAYER metal3 ;
  RECT 1833.120 0.000 1836.660 1.120 ;
  LAYER metal2 ;
  RECT 1833.120 0.000 1836.660 1.120 ;
  LAYER metal1 ;
  RECT 1833.120 0.000 1836.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1803.980 0.000 1807.520 1.120 ;
  LAYER metal4 ;
  RECT 1803.980 0.000 1807.520 1.120 ;
  LAYER metal3 ;
  RECT 1803.980 0.000 1807.520 1.120 ;
  LAYER metal2 ;
  RECT 1803.980 0.000 1807.520 1.120 ;
  LAYER metal1 ;
  RECT 1803.980 0.000 1807.520 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1779.800 0.000 1783.340 1.120 ;
  LAYER metal4 ;
  RECT 1779.800 0.000 1783.340 1.120 ;
  LAYER metal3 ;
  RECT 1779.800 0.000 1783.340 1.120 ;
  LAYER metal2 ;
  RECT 1779.800 0.000 1783.340 1.120 ;
  LAYER metal1 ;
  RECT 1779.800 0.000 1783.340 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1756.860 0.000 1760.400 1.120 ;
  LAYER metal4 ;
  RECT 1756.860 0.000 1760.400 1.120 ;
  LAYER metal3 ;
  RECT 1756.860 0.000 1760.400 1.120 ;
  LAYER metal2 ;
  RECT 1756.860 0.000 1760.400 1.120 ;
  LAYER metal1 ;
  RECT 1756.860 0.000 1760.400 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1748.180 0.000 1751.720 1.120 ;
  LAYER metal4 ;
  RECT 1748.180 0.000 1751.720 1.120 ;
  LAYER metal3 ;
  RECT 1748.180 0.000 1751.720 1.120 ;
  LAYER metal2 ;
  RECT 1748.180 0.000 1751.720 1.120 ;
  LAYER metal1 ;
  RECT 1748.180 0.000 1751.720 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1685.560 0.000 1689.100 1.120 ;
  LAYER metal4 ;
  RECT 1685.560 0.000 1689.100 1.120 ;
  LAYER metal3 ;
  RECT 1685.560 0.000 1689.100 1.120 ;
  LAYER metal2 ;
  RECT 1685.560 0.000 1689.100 1.120 ;
  LAYER metal1 ;
  RECT 1685.560 0.000 1689.100 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1672.540 0.000 1676.080 1.120 ;
  LAYER metal4 ;
  RECT 1672.540 0.000 1676.080 1.120 ;
  LAYER metal3 ;
  RECT 1672.540 0.000 1676.080 1.120 ;
  LAYER metal2 ;
  RECT 1672.540 0.000 1676.080 1.120 ;
  LAYER metal1 ;
  RECT 1672.540 0.000 1676.080 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1658.900 0.000 1662.440 1.120 ;
  LAYER metal4 ;
  RECT 1658.900 0.000 1662.440 1.120 ;
  LAYER metal3 ;
  RECT 1658.900 0.000 1662.440 1.120 ;
  LAYER metal2 ;
  RECT 1658.900 0.000 1662.440 1.120 ;
  LAYER metal1 ;
  RECT 1658.900 0.000 1662.440 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1645.260 0.000 1648.800 1.120 ;
  LAYER metal4 ;
  RECT 1645.260 0.000 1648.800 1.120 ;
  LAYER metal3 ;
  RECT 1645.260 0.000 1648.800 1.120 ;
  LAYER metal2 ;
  RECT 1645.260 0.000 1648.800 1.120 ;
  LAYER metal1 ;
  RECT 1645.260 0.000 1648.800 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1632.240 0.000 1635.780 1.120 ;
  LAYER metal4 ;
  RECT 1632.240 0.000 1635.780 1.120 ;
  LAYER metal3 ;
  RECT 1632.240 0.000 1635.780 1.120 ;
  LAYER metal2 ;
  RECT 1632.240 0.000 1635.780 1.120 ;
  LAYER metal1 ;
  RECT 1632.240 0.000 1635.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1618.600 0.000 1622.140 1.120 ;
  LAYER metal4 ;
  RECT 1618.600 0.000 1622.140 1.120 ;
  LAYER metal3 ;
  RECT 1618.600 0.000 1622.140 1.120 ;
  LAYER metal2 ;
  RECT 1618.600 0.000 1622.140 1.120 ;
  LAYER metal1 ;
  RECT 1618.600 0.000 1622.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1551.640 0.000 1555.180 1.120 ;
  LAYER metal4 ;
  RECT 1551.640 0.000 1555.180 1.120 ;
  LAYER metal3 ;
  RECT 1551.640 0.000 1555.180 1.120 ;
  LAYER metal2 ;
  RECT 1551.640 0.000 1555.180 1.120 ;
  LAYER metal1 ;
  RECT 1551.640 0.000 1555.180 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1538.000 0.000 1541.540 1.120 ;
  LAYER metal4 ;
  RECT 1538.000 0.000 1541.540 1.120 ;
  LAYER metal3 ;
  RECT 1538.000 0.000 1541.540 1.120 ;
  LAYER metal2 ;
  RECT 1538.000 0.000 1541.540 1.120 ;
  LAYER metal1 ;
  RECT 1538.000 0.000 1541.540 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1524.360 0.000 1527.900 1.120 ;
  LAYER metal4 ;
  RECT 1524.360 0.000 1527.900 1.120 ;
  LAYER metal3 ;
  RECT 1524.360 0.000 1527.900 1.120 ;
  LAYER metal2 ;
  RECT 1524.360 0.000 1527.900 1.120 ;
  LAYER metal1 ;
  RECT 1524.360 0.000 1527.900 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1511.340 0.000 1514.880 1.120 ;
  LAYER metal4 ;
  RECT 1511.340 0.000 1514.880 1.120 ;
  LAYER metal3 ;
  RECT 1511.340 0.000 1514.880 1.120 ;
  LAYER metal2 ;
  RECT 1511.340 0.000 1514.880 1.120 ;
  LAYER metal1 ;
  RECT 1511.340 0.000 1514.880 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1497.700 0.000 1501.240 1.120 ;
  LAYER metal4 ;
  RECT 1497.700 0.000 1501.240 1.120 ;
  LAYER metal3 ;
  RECT 1497.700 0.000 1501.240 1.120 ;
  LAYER metal2 ;
  RECT 1497.700 0.000 1501.240 1.120 ;
  LAYER metal1 ;
  RECT 1497.700 0.000 1501.240 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1484.060 0.000 1487.600 1.120 ;
  LAYER metal4 ;
  RECT 1484.060 0.000 1487.600 1.120 ;
  LAYER metal3 ;
  RECT 1484.060 0.000 1487.600 1.120 ;
  LAYER metal2 ;
  RECT 1484.060 0.000 1487.600 1.120 ;
  LAYER metal1 ;
  RECT 1484.060 0.000 1487.600 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1417.100 0.000 1420.640 1.120 ;
  LAYER metal4 ;
  RECT 1417.100 0.000 1420.640 1.120 ;
  LAYER metal3 ;
  RECT 1417.100 0.000 1420.640 1.120 ;
  LAYER metal2 ;
  RECT 1417.100 0.000 1420.640 1.120 ;
  LAYER metal1 ;
  RECT 1417.100 0.000 1420.640 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1403.460 0.000 1407.000 1.120 ;
  LAYER metal4 ;
  RECT 1403.460 0.000 1407.000 1.120 ;
  LAYER metal3 ;
  RECT 1403.460 0.000 1407.000 1.120 ;
  LAYER metal2 ;
  RECT 1403.460 0.000 1407.000 1.120 ;
  LAYER metal1 ;
  RECT 1403.460 0.000 1407.000 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1390.440 0.000 1393.980 1.120 ;
  LAYER metal4 ;
  RECT 1390.440 0.000 1393.980 1.120 ;
  LAYER metal3 ;
  RECT 1390.440 0.000 1393.980 1.120 ;
  LAYER metal2 ;
  RECT 1390.440 0.000 1393.980 1.120 ;
  LAYER metal1 ;
  RECT 1390.440 0.000 1393.980 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1376.800 0.000 1380.340 1.120 ;
  LAYER metal4 ;
  RECT 1376.800 0.000 1380.340 1.120 ;
  LAYER metal3 ;
  RECT 1376.800 0.000 1380.340 1.120 ;
  LAYER metal2 ;
  RECT 1376.800 0.000 1380.340 1.120 ;
  LAYER metal1 ;
  RECT 1376.800 0.000 1380.340 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1363.160 0.000 1366.700 1.120 ;
  LAYER metal4 ;
  RECT 1363.160 0.000 1366.700 1.120 ;
  LAYER metal3 ;
  RECT 1363.160 0.000 1366.700 1.120 ;
  LAYER metal2 ;
  RECT 1363.160 0.000 1366.700 1.120 ;
  LAYER metal1 ;
  RECT 1363.160 0.000 1366.700 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1350.140 0.000 1353.680 1.120 ;
  LAYER metal4 ;
  RECT 1350.140 0.000 1353.680 1.120 ;
  LAYER metal3 ;
  RECT 1350.140 0.000 1353.680 1.120 ;
  LAYER metal2 ;
  RECT 1350.140 0.000 1353.680 1.120 ;
  LAYER metal1 ;
  RECT 1350.140 0.000 1353.680 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1282.560 0.000 1286.100 1.120 ;
  LAYER metal4 ;
  RECT 1282.560 0.000 1286.100 1.120 ;
  LAYER metal3 ;
  RECT 1282.560 0.000 1286.100 1.120 ;
  LAYER metal2 ;
  RECT 1282.560 0.000 1286.100 1.120 ;
  LAYER metal1 ;
  RECT 1282.560 0.000 1286.100 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1268.920 0.000 1272.460 1.120 ;
  LAYER metal4 ;
  RECT 1268.920 0.000 1272.460 1.120 ;
  LAYER metal3 ;
  RECT 1268.920 0.000 1272.460 1.120 ;
  LAYER metal2 ;
  RECT 1268.920 0.000 1272.460 1.120 ;
  LAYER metal1 ;
  RECT 1268.920 0.000 1272.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1255.900 0.000 1259.440 1.120 ;
  LAYER metal4 ;
  RECT 1255.900 0.000 1259.440 1.120 ;
  LAYER metal3 ;
  RECT 1255.900 0.000 1259.440 1.120 ;
  LAYER metal2 ;
  RECT 1255.900 0.000 1259.440 1.120 ;
  LAYER metal1 ;
  RECT 1255.900 0.000 1259.440 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1242.260 0.000 1245.800 1.120 ;
  LAYER metal4 ;
  RECT 1242.260 0.000 1245.800 1.120 ;
  LAYER metal3 ;
  RECT 1242.260 0.000 1245.800 1.120 ;
  LAYER metal2 ;
  RECT 1242.260 0.000 1245.800 1.120 ;
  LAYER metal1 ;
  RECT 1242.260 0.000 1245.800 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1228.620 0.000 1232.160 1.120 ;
  LAYER metal4 ;
  RECT 1228.620 0.000 1232.160 1.120 ;
  LAYER metal3 ;
  RECT 1228.620 0.000 1232.160 1.120 ;
  LAYER metal2 ;
  RECT 1228.620 0.000 1232.160 1.120 ;
  LAYER metal1 ;
  RECT 1228.620 0.000 1232.160 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1215.600 0.000 1219.140 1.120 ;
  LAYER metal4 ;
  RECT 1215.600 0.000 1219.140 1.120 ;
  LAYER metal3 ;
  RECT 1215.600 0.000 1219.140 1.120 ;
  LAYER metal2 ;
  RECT 1215.600 0.000 1219.140 1.120 ;
  LAYER metal1 ;
  RECT 1215.600 0.000 1219.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1148.020 0.000 1151.560 1.120 ;
  LAYER metal4 ;
  RECT 1148.020 0.000 1151.560 1.120 ;
  LAYER metal3 ;
  RECT 1148.020 0.000 1151.560 1.120 ;
  LAYER metal2 ;
  RECT 1148.020 0.000 1151.560 1.120 ;
  LAYER metal1 ;
  RECT 1148.020 0.000 1151.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1135.000 0.000 1138.540 1.120 ;
  LAYER metal4 ;
  RECT 1135.000 0.000 1138.540 1.120 ;
  LAYER metal3 ;
  RECT 1135.000 0.000 1138.540 1.120 ;
  LAYER metal2 ;
  RECT 1135.000 0.000 1138.540 1.120 ;
  LAYER metal1 ;
  RECT 1135.000 0.000 1138.540 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1121.360 0.000 1124.900 1.120 ;
  LAYER metal4 ;
  RECT 1121.360 0.000 1124.900 1.120 ;
  LAYER metal3 ;
  RECT 1121.360 0.000 1124.900 1.120 ;
  LAYER metal2 ;
  RECT 1121.360 0.000 1124.900 1.120 ;
  LAYER metal1 ;
  RECT 1121.360 0.000 1124.900 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1107.720 0.000 1111.260 1.120 ;
  LAYER metal4 ;
  RECT 1107.720 0.000 1111.260 1.120 ;
  LAYER metal3 ;
  RECT 1107.720 0.000 1111.260 1.120 ;
  LAYER metal2 ;
  RECT 1107.720 0.000 1111.260 1.120 ;
  LAYER metal1 ;
  RECT 1107.720 0.000 1111.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1094.700 0.000 1098.240 1.120 ;
  LAYER metal4 ;
  RECT 1094.700 0.000 1098.240 1.120 ;
  LAYER metal3 ;
  RECT 1094.700 0.000 1098.240 1.120 ;
  LAYER metal2 ;
  RECT 1094.700 0.000 1098.240 1.120 ;
  LAYER metal1 ;
  RECT 1094.700 0.000 1098.240 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1081.060 0.000 1084.600 1.120 ;
  LAYER metal4 ;
  RECT 1081.060 0.000 1084.600 1.120 ;
  LAYER metal3 ;
  RECT 1081.060 0.000 1084.600 1.120 ;
  LAYER metal2 ;
  RECT 1081.060 0.000 1084.600 1.120 ;
  LAYER metal1 ;
  RECT 1081.060 0.000 1084.600 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1014.100 0.000 1017.640 1.120 ;
  LAYER metal4 ;
  RECT 1014.100 0.000 1017.640 1.120 ;
  LAYER metal3 ;
  RECT 1014.100 0.000 1017.640 1.120 ;
  LAYER metal2 ;
  RECT 1014.100 0.000 1017.640 1.120 ;
  LAYER metal1 ;
  RECT 1014.100 0.000 1017.640 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1000.460 0.000 1004.000 1.120 ;
  LAYER metal4 ;
  RECT 1000.460 0.000 1004.000 1.120 ;
  LAYER metal3 ;
  RECT 1000.460 0.000 1004.000 1.120 ;
  LAYER metal2 ;
  RECT 1000.460 0.000 1004.000 1.120 ;
  LAYER metal1 ;
  RECT 1000.460 0.000 1004.000 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 986.820 0.000 990.360 1.120 ;
  LAYER metal4 ;
  RECT 986.820 0.000 990.360 1.120 ;
  LAYER metal3 ;
  RECT 986.820 0.000 990.360 1.120 ;
  LAYER metal2 ;
  RECT 986.820 0.000 990.360 1.120 ;
  LAYER metal1 ;
  RECT 986.820 0.000 990.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 973.800 0.000 977.340 1.120 ;
  LAYER metal4 ;
  RECT 973.800 0.000 977.340 1.120 ;
  LAYER metal3 ;
  RECT 973.800 0.000 977.340 1.120 ;
  LAYER metal2 ;
  RECT 973.800 0.000 977.340 1.120 ;
  LAYER metal1 ;
  RECT 973.800 0.000 977.340 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 960.160 0.000 963.700 1.120 ;
  LAYER metal4 ;
  RECT 960.160 0.000 963.700 1.120 ;
  LAYER metal3 ;
  RECT 960.160 0.000 963.700 1.120 ;
  LAYER metal2 ;
  RECT 960.160 0.000 963.700 1.120 ;
  LAYER metal1 ;
  RECT 960.160 0.000 963.700 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 946.520 0.000 950.060 1.120 ;
  LAYER metal4 ;
  RECT 946.520 0.000 950.060 1.120 ;
  LAYER metal3 ;
  RECT 946.520 0.000 950.060 1.120 ;
  LAYER metal2 ;
  RECT 946.520 0.000 950.060 1.120 ;
  LAYER metal1 ;
  RECT 946.520 0.000 950.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 879.560 0.000 883.100 1.120 ;
  LAYER metal4 ;
  RECT 879.560 0.000 883.100 1.120 ;
  LAYER metal3 ;
  RECT 879.560 0.000 883.100 1.120 ;
  LAYER metal2 ;
  RECT 879.560 0.000 883.100 1.120 ;
  LAYER metal1 ;
  RECT 879.560 0.000 883.100 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 865.920 0.000 869.460 1.120 ;
  LAYER metal4 ;
  RECT 865.920 0.000 869.460 1.120 ;
  LAYER metal3 ;
  RECT 865.920 0.000 869.460 1.120 ;
  LAYER metal2 ;
  RECT 865.920 0.000 869.460 1.120 ;
  LAYER metal1 ;
  RECT 865.920 0.000 869.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 852.280 0.000 855.820 1.120 ;
  LAYER metal4 ;
  RECT 852.280 0.000 855.820 1.120 ;
  LAYER metal3 ;
  RECT 852.280 0.000 855.820 1.120 ;
  LAYER metal2 ;
  RECT 852.280 0.000 855.820 1.120 ;
  LAYER metal1 ;
  RECT 852.280 0.000 855.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 839.260 0.000 842.800 1.120 ;
  LAYER metal4 ;
  RECT 839.260 0.000 842.800 1.120 ;
  LAYER metal3 ;
  RECT 839.260 0.000 842.800 1.120 ;
  LAYER metal2 ;
  RECT 839.260 0.000 842.800 1.120 ;
  LAYER metal1 ;
  RECT 839.260 0.000 842.800 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 825.620 0.000 829.160 1.120 ;
  LAYER metal4 ;
  RECT 825.620 0.000 829.160 1.120 ;
  LAYER metal3 ;
  RECT 825.620 0.000 829.160 1.120 ;
  LAYER metal2 ;
  RECT 825.620 0.000 829.160 1.120 ;
  LAYER metal1 ;
  RECT 825.620 0.000 829.160 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 811.980 0.000 815.520 1.120 ;
  LAYER metal4 ;
  RECT 811.980 0.000 815.520 1.120 ;
  LAYER metal3 ;
  RECT 811.980 0.000 815.520 1.120 ;
  LAYER metal2 ;
  RECT 811.980 0.000 815.520 1.120 ;
  LAYER metal1 ;
  RECT 811.980 0.000 815.520 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 745.020 0.000 748.560 1.120 ;
  LAYER metal4 ;
  RECT 745.020 0.000 748.560 1.120 ;
  LAYER metal3 ;
  RECT 745.020 0.000 748.560 1.120 ;
  LAYER metal2 ;
  RECT 745.020 0.000 748.560 1.120 ;
  LAYER metal1 ;
  RECT 745.020 0.000 748.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 731.380 0.000 734.920 1.120 ;
  LAYER metal4 ;
  RECT 731.380 0.000 734.920 1.120 ;
  LAYER metal3 ;
  RECT 731.380 0.000 734.920 1.120 ;
  LAYER metal2 ;
  RECT 731.380 0.000 734.920 1.120 ;
  LAYER metal1 ;
  RECT 731.380 0.000 734.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 718.360 0.000 721.900 1.120 ;
  LAYER metal4 ;
  RECT 718.360 0.000 721.900 1.120 ;
  LAYER metal3 ;
  RECT 718.360 0.000 721.900 1.120 ;
  LAYER metal2 ;
  RECT 718.360 0.000 721.900 1.120 ;
  LAYER metal1 ;
  RECT 718.360 0.000 721.900 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 704.720 0.000 708.260 1.120 ;
  LAYER metal4 ;
  RECT 704.720 0.000 708.260 1.120 ;
  LAYER metal3 ;
  RECT 704.720 0.000 708.260 1.120 ;
  LAYER metal2 ;
  RECT 704.720 0.000 708.260 1.120 ;
  LAYER metal1 ;
  RECT 704.720 0.000 708.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 691.080 0.000 694.620 1.120 ;
  LAYER metal4 ;
  RECT 691.080 0.000 694.620 1.120 ;
  LAYER metal3 ;
  RECT 691.080 0.000 694.620 1.120 ;
  LAYER metal2 ;
  RECT 691.080 0.000 694.620 1.120 ;
  LAYER metal1 ;
  RECT 691.080 0.000 694.620 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 678.060 0.000 681.600 1.120 ;
  LAYER metal4 ;
  RECT 678.060 0.000 681.600 1.120 ;
  LAYER metal3 ;
  RECT 678.060 0.000 681.600 1.120 ;
  LAYER metal2 ;
  RECT 678.060 0.000 681.600 1.120 ;
  LAYER metal1 ;
  RECT 678.060 0.000 681.600 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 610.480 0.000 614.020 1.120 ;
  LAYER metal4 ;
  RECT 610.480 0.000 614.020 1.120 ;
  LAYER metal3 ;
  RECT 610.480 0.000 614.020 1.120 ;
  LAYER metal2 ;
  RECT 610.480 0.000 614.020 1.120 ;
  LAYER metal1 ;
  RECT 610.480 0.000 614.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 597.460 0.000 601.000 1.120 ;
  LAYER metal4 ;
  RECT 597.460 0.000 601.000 1.120 ;
  LAYER metal3 ;
  RECT 597.460 0.000 601.000 1.120 ;
  LAYER metal2 ;
  RECT 597.460 0.000 601.000 1.120 ;
  LAYER metal1 ;
  RECT 597.460 0.000 601.000 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 583.820 0.000 587.360 1.120 ;
  LAYER metal4 ;
  RECT 583.820 0.000 587.360 1.120 ;
  LAYER metal3 ;
  RECT 583.820 0.000 587.360 1.120 ;
  LAYER metal2 ;
  RECT 583.820 0.000 587.360 1.120 ;
  LAYER metal1 ;
  RECT 583.820 0.000 587.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 570.180 0.000 573.720 1.120 ;
  LAYER metal4 ;
  RECT 570.180 0.000 573.720 1.120 ;
  LAYER metal3 ;
  RECT 570.180 0.000 573.720 1.120 ;
  LAYER metal2 ;
  RECT 570.180 0.000 573.720 1.120 ;
  LAYER metal1 ;
  RECT 570.180 0.000 573.720 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 557.160 0.000 560.700 1.120 ;
  LAYER metal4 ;
  RECT 557.160 0.000 560.700 1.120 ;
  LAYER metal3 ;
  RECT 557.160 0.000 560.700 1.120 ;
  LAYER metal2 ;
  RECT 557.160 0.000 560.700 1.120 ;
  LAYER metal1 ;
  RECT 557.160 0.000 560.700 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 543.520 0.000 547.060 1.120 ;
  LAYER metal4 ;
  RECT 543.520 0.000 547.060 1.120 ;
  LAYER metal3 ;
  RECT 543.520 0.000 547.060 1.120 ;
  LAYER metal2 ;
  RECT 543.520 0.000 547.060 1.120 ;
  LAYER metal1 ;
  RECT 543.520 0.000 547.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 475.940 0.000 479.480 1.120 ;
  LAYER metal4 ;
  RECT 475.940 0.000 479.480 1.120 ;
  LAYER metal3 ;
  RECT 475.940 0.000 479.480 1.120 ;
  LAYER metal2 ;
  RECT 475.940 0.000 479.480 1.120 ;
  LAYER metal1 ;
  RECT 475.940 0.000 479.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 462.920 0.000 466.460 1.120 ;
  LAYER metal4 ;
  RECT 462.920 0.000 466.460 1.120 ;
  LAYER metal3 ;
  RECT 462.920 0.000 466.460 1.120 ;
  LAYER metal2 ;
  RECT 462.920 0.000 466.460 1.120 ;
  LAYER metal1 ;
  RECT 462.920 0.000 466.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 449.280 0.000 452.820 1.120 ;
  LAYER metal4 ;
  RECT 449.280 0.000 452.820 1.120 ;
  LAYER metal3 ;
  RECT 449.280 0.000 452.820 1.120 ;
  LAYER metal2 ;
  RECT 449.280 0.000 452.820 1.120 ;
  LAYER metal1 ;
  RECT 449.280 0.000 452.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 435.640 0.000 439.180 1.120 ;
  LAYER metal4 ;
  RECT 435.640 0.000 439.180 1.120 ;
  LAYER metal3 ;
  RECT 435.640 0.000 439.180 1.120 ;
  LAYER metal2 ;
  RECT 435.640 0.000 439.180 1.120 ;
  LAYER metal1 ;
  RECT 435.640 0.000 439.180 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 422.620 0.000 426.160 1.120 ;
  LAYER metal4 ;
  RECT 422.620 0.000 426.160 1.120 ;
  LAYER metal3 ;
  RECT 422.620 0.000 426.160 1.120 ;
  LAYER metal2 ;
  RECT 422.620 0.000 426.160 1.120 ;
  LAYER metal1 ;
  RECT 422.620 0.000 426.160 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 408.980 0.000 412.520 1.120 ;
  LAYER metal4 ;
  RECT 408.980 0.000 412.520 1.120 ;
  LAYER metal3 ;
  RECT 408.980 0.000 412.520 1.120 ;
  LAYER metal2 ;
  RECT 408.980 0.000 412.520 1.120 ;
  LAYER metal1 ;
  RECT 408.980 0.000 412.520 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 342.020 0.000 345.560 1.120 ;
  LAYER metal4 ;
  RECT 342.020 0.000 345.560 1.120 ;
  LAYER metal3 ;
  RECT 342.020 0.000 345.560 1.120 ;
  LAYER metal2 ;
  RECT 342.020 0.000 345.560 1.120 ;
  LAYER metal1 ;
  RECT 342.020 0.000 345.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 328.380 0.000 331.920 1.120 ;
  LAYER metal4 ;
  RECT 328.380 0.000 331.920 1.120 ;
  LAYER metal3 ;
  RECT 328.380 0.000 331.920 1.120 ;
  LAYER metal2 ;
  RECT 328.380 0.000 331.920 1.120 ;
  LAYER metal1 ;
  RECT 328.380 0.000 331.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 314.740 0.000 318.280 1.120 ;
  LAYER metal4 ;
  RECT 314.740 0.000 318.280 1.120 ;
  LAYER metal3 ;
  RECT 314.740 0.000 318.280 1.120 ;
  LAYER metal2 ;
  RECT 314.740 0.000 318.280 1.120 ;
  LAYER metal1 ;
  RECT 314.740 0.000 318.280 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 301.720 0.000 305.260 1.120 ;
  LAYER metal4 ;
  RECT 301.720 0.000 305.260 1.120 ;
  LAYER metal3 ;
  RECT 301.720 0.000 305.260 1.120 ;
  LAYER metal2 ;
  RECT 301.720 0.000 305.260 1.120 ;
  LAYER metal1 ;
  RECT 301.720 0.000 305.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 288.080 0.000 291.620 1.120 ;
  LAYER metal4 ;
  RECT 288.080 0.000 291.620 1.120 ;
  LAYER metal3 ;
  RECT 288.080 0.000 291.620 1.120 ;
  LAYER metal2 ;
  RECT 288.080 0.000 291.620 1.120 ;
  LAYER metal1 ;
  RECT 288.080 0.000 291.620 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 274.440 0.000 277.980 1.120 ;
  LAYER metal4 ;
  RECT 274.440 0.000 277.980 1.120 ;
  LAYER metal3 ;
  RECT 274.440 0.000 277.980 1.120 ;
  LAYER metal2 ;
  RECT 274.440 0.000 277.980 1.120 ;
  LAYER metal1 ;
  RECT 274.440 0.000 277.980 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 207.480 0.000 211.020 1.120 ;
  LAYER metal4 ;
  RECT 207.480 0.000 211.020 1.120 ;
  LAYER metal3 ;
  RECT 207.480 0.000 211.020 1.120 ;
  LAYER metal2 ;
  RECT 207.480 0.000 211.020 1.120 ;
  LAYER metal1 ;
  RECT 207.480 0.000 211.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 193.840 0.000 197.380 1.120 ;
  LAYER metal4 ;
  RECT 193.840 0.000 197.380 1.120 ;
  LAYER metal3 ;
  RECT 193.840 0.000 197.380 1.120 ;
  LAYER metal2 ;
  RECT 193.840 0.000 197.380 1.120 ;
  LAYER metal1 ;
  RECT 193.840 0.000 197.380 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 180.820 0.000 184.360 1.120 ;
  LAYER metal4 ;
  RECT 180.820 0.000 184.360 1.120 ;
  LAYER metal3 ;
  RECT 180.820 0.000 184.360 1.120 ;
  LAYER metal2 ;
  RECT 180.820 0.000 184.360 1.120 ;
  LAYER metal1 ;
  RECT 180.820 0.000 184.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 167.180 0.000 170.720 1.120 ;
  LAYER metal4 ;
  RECT 167.180 0.000 170.720 1.120 ;
  LAYER metal3 ;
  RECT 167.180 0.000 170.720 1.120 ;
  LAYER metal2 ;
  RECT 167.180 0.000 170.720 1.120 ;
  LAYER metal1 ;
  RECT 167.180 0.000 170.720 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 153.540 0.000 157.080 1.120 ;
  LAYER metal4 ;
  RECT 153.540 0.000 157.080 1.120 ;
  LAYER metal3 ;
  RECT 153.540 0.000 157.080 1.120 ;
  LAYER metal2 ;
  RECT 153.540 0.000 157.080 1.120 ;
  LAYER metal1 ;
  RECT 153.540 0.000 157.080 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 140.520 0.000 144.060 1.120 ;
  LAYER metal4 ;
  RECT 140.520 0.000 144.060 1.120 ;
  LAYER metal3 ;
  RECT 140.520 0.000 144.060 1.120 ;
  LAYER metal2 ;
  RECT 140.520 0.000 144.060 1.120 ;
  LAYER metal1 ;
  RECT 140.520 0.000 144.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 72.940 0.000 76.480 1.120 ;
  LAYER metal4 ;
  RECT 72.940 0.000 76.480 1.120 ;
  LAYER metal3 ;
  RECT 72.940 0.000 76.480 1.120 ;
  LAYER metal2 ;
  RECT 72.940 0.000 76.480 1.120 ;
  LAYER metal1 ;
  RECT 72.940 0.000 76.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 59.300 0.000 62.840 1.120 ;
  LAYER metal4 ;
  RECT 59.300 0.000 62.840 1.120 ;
  LAYER metal3 ;
  RECT 59.300 0.000 62.840 1.120 ;
  LAYER metal2 ;
  RECT 59.300 0.000 62.840 1.120 ;
  LAYER metal1 ;
  RECT 59.300 0.000 62.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 46.280 0.000 49.820 1.120 ;
  LAYER metal4 ;
  RECT 46.280 0.000 49.820 1.120 ;
  LAYER metal3 ;
  RECT 46.280 0.000 49.820 1.120 ;
  LAYER metal2 ;
  RECT 46.280 0.000 49.820 1.120 ;
  LAYER metal1 ;
  RECT 46.280 0.000 49.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 32.640 0.000 36.180 1.120 ;
  LAYER metal4 ;
  RECT 32.640 0.000 36.180 1.120 ;
  LAYER metal3 ;
  RECT 32.640 0.000 36.180 1.120 ;
  LAYER metal2 ;
  RECT 32.640 0.000 36.180 1.120 ;
  LAYER metal1 ;
  RECT 32.640 0.000 36.180 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 19.000 0.000 22.540 1.120 ;
  LAYER metal4 ;
  RECT 19.000 0.000 22.540 1.120 ;
  LAYER metal3 ;
  RECT 19.000 0.000 22.540 1.120 ;
  LAYER metal2 ;
  RECT 19.000 0.000 22.540 1.120 ;
  LAYER metal1 ;
  RECT 19.000 0.000 22.540 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 7.220 0.000 10.760 1.120 ;
  LAYER metal4 ;
  RECT 7.220 0.000 10.760 1.120 ;
  LAYER metal3 ;
  RECT 7.220 0.000 10.760 1.120 ;
  LAYER metal2 ;
  RECT 7.220 0.000 10.760 1.120 ;
  LAYER metal1 ;
  RECT 7.220 0.000 10.760 1.120 ;
 END
END VCC
PIN DIB127
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3573.120 500.640 3574.240 501.760 ;
  LAYER metal4 ;
  RECT 3573.120 500.640 3574.240 501.760 ;
  LAYER metal3 ;
  RECT 3573.120 500.640 3574.240 501.760 ;
  LAYER metal2 ;
  RECT 3573.120 500.640 3574.240 501.760 ;
  LAYER metal1 ;
  RECT 3573.120 500.640 3574.240 501.760 ;
 END
END DIB127
PIN DOB127
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3559.480 500.640 3560.600 501.760 ;
  LAYER metal4 ;
  RECT 3559.480 500.640 3560.600 501.760 ;
  LAYER metal3 ;
  RECT 3559.480 500.640 3560.600 501.760 ;
  LAYER metal2 ;
  RECT 3559.480 500.640 3560.600 501.760 ;
  LAYER metal1 ;
  RECT 3559.480 500.640 3560.600 501.760 ;
 END
END DOB127
PIN DIB126
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3546.460 500.640 3547.580 501.760 ;
  LAYER metal4 ;
  RECT 3546.460 500.640 3547.580 501.760 ;
  LAYER metal3 ;
  RECT 3546.460 500.640 3547.580 501.760 ;
  LAYER metal2 ;
  RECT 3546.460 500.640 3547.580 501.760 ;
  LAYER metal1 ;
  RECT 3546.460 500.640 3547.580 501.760 ;
 END
END DIB126
PIN DOB126
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3532.820 500.640 3533.940 501.760 ;
  LAYER metal4 ;
  RECT 3532.820 500.640 3533.940 501.760 ;
  LAYER metal3 ;
  RECT 3532.820 500.640 3533.940 501.760 ;
  LAYER metal2 ;
  RECT 3532.820 500.640 3533.940 501.760 ;
  LAYER metal1 ;
  RECT 3532.820 500.640 3533.940 501.760 ;
 END
END DOB126
PIN DIB125
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3519.180 500.640 3520.300 501.760 ;
  LAYER metal4 ;
  RECT 3519.180 500.640 3520.300 501.760 ;
  LAYER metal3 ;
  RECT 3519.180 500.640 3520.300 501.760 ;
  LAYER metal2 ;
  RECT 3519.180 500.640 3520.300 501.760 ;
  LAYER metal1 ;
  RECT 3519.180 500.640 3520.300 501.760 ;
 END
END DIB125
PIN DOB125
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3506.160 500.640 3507.280 501.760 ;
  LAYER metal4 ;
  RECT 3506.160 500.640 3507.280 501.760 ;
  LAYER metal3 ;
  RECT 3506.160 500.640 3507.280 501.760 ;
  LAYER metal2 ;
  RECT 3506.160 500.640 3507.280 501.760 ;
  LAYER metal1 ;
  RECT 3506.160 500.640 3507.280 501.760 ;
 END
END DOB125
PIN DIB124
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3492.520 500.640 3493.640 501.760 ;
  LAYER metal4 ;
  RECT 3492.520 500.640 3493.640 501.760 ;
  LAYER metal3 ;
  RECT 3492.520 500.640 3493.640 501.760 ;
  LAYER metal2 ;
  RECT 3492.520 500.640 3493.640 501.760 ;
  LAYER metal1 ;
  RECT 3492.520 500.640 3493.640 501.760 ;
 END
END DIB124
PIN DOB124
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3478.880 500.640 3480.000 501.760 ;
  LAYER metal4 ;
  RECT 3478.880 500.640 3480.000 501.760 ;
  LAYER metal3 ;
  RECT 3478.880 500.640 3480.000 501.760 ;
  LAYER metal2 ;
  RECT 3478.880 500.640 3480.000 501.760 ;
  LAYER metal1 ;
  RECT 3478.880 500.640 3480.000 501.760 ;
 END
END DOB124
PIN DIB123
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3465.860 500.640 3466.980 501.760 ;
  LAYER metal4 ;
  RECT 3465.860 500.640 3466.980 501.760 ;
  LAYER metal3 ;
  RECT 3465.860 500.640 3466.980 501.760 ;
  LAYER metal2 ;
  RECT 3465.860 500.640 3466.980 501.760 ;
  LAYER metal1 ;
  RECT 3465.860 500.640 3466.980 501.760 ;
 END
END DIB123
PIN DOB123
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3452.220 500.640 3453.340 501.760 ;
  LAYER metal4 ;
  RECT 3452.220 500.640 3453.340 501.760 ;
  LAYER metal3 ;
  RECT 3452.220 500.640 3453.340 501.760 ;
  LAYER metal2 ;
  RECT 3452.220 500.640 3453.340 501.760 ;
  LAYER metal1 ;
  RECT 3452.220 500.640 3453.340 501.760 ;
 END
END DOB123
PIN DIB122
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3438.580 500.640 3439.700 501.760 ;
  LAYER metal4 ;
  RECT 3438.580 500.640 3439.700 501.760 ;
  LAYER metal3 ;
  RECT 3438.580 500.640 3439.700 501.760 ;
  LAYER metal2 ;
  RECT 3438.580 500.640 3439.700 501.760 ;
  LAYER metal1 ;
  RECT 3438.580 500.640 3439.700 501.760 ;
 END
END DIB122
PIN DOB122
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3425.560 500.640 3426.680 501.760 ;
  LAYER metal4 ;
  RECT 3425.560 500.640 3426.680 501.760 ;
  LAYER metal3 ;
  RECT 3425.560 500.640 3426.680 501.760 ;
  LAYER metal2 ;
  RECT 3425.560 500.640 3426.680 501.760 ;
  LAYER metal1 ;
  RECT 3425.560 500.640 3426.680 501.760 ;
 END
END DOB122
PIN DIB121
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3411.920 500.640 3413.040 501.760 ;
  LAYER metal4 ;
  RECT 3411.920 500.640 3413.040 501.760 ;
  LAYER metal3 ;
  RECT 3411.920 500.640 3413.040 501.760 ;
  LAYER metal2 ;
  RECT 3411.920 500.640 3413.040 501.760 ;
  LAYER metal1 ;
  RECT 3411.920 500.640 3413.040 501.760 ;
 END
END DIB121
PIN DOB121
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3398.280 500.640 3399.400 501.760 ;
  LAYER metal4 ;
  RECT 3398.280 500.640 3399.400 501.760 ;
  LAYER metal3 ;
  RECT 3398.280 500.640 3399.400 501.760 ;
  LAYER metal2 ;
  RECT 3398.280 500.640 3399.400 501.760 ;
  LAYER metal1 ;
  RECT 3398.280 500.640 3399.400 501.760 ;
 END
END DOB121
PIN DIB120
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3385.260 500.640 3386.380 501.760 ;
  LAYER metal4 ;
  RECT 3385.260 500.640 3386.380 501.760 ;
  LAYER metal3 ;
  RECT 3385.260 500.640 3386.380 501.760 ;
  LAYER metal2 ;
  RECT 3385.260 500.640 3386.380 501.760 ;
  LAYER metal1 ;
  RECT 3385.260 500.640 3386.380 501.760 ;
 END
END DIB120
PIN DOB120
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3371.620 500.640 3372.740 501.760 ;
  LAYER metal4 ;
  RECT 3371.620 500.640 3372.740 501.760 ;
  LAYER metal3 ;
  RECT 3371.620 500.640 3372.740 501.760 ;
  LAYER metal2 ;
  RECT 3371.620 500.640 3372.740 501.760 ;
  LAYER metal1 ;
  RECT 3371.620 500.640 3372.740 501.760 ;
 END
END DOB120
PIN DIB119
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3357.980 500.640 3359.100 501.760 ;
  LAYER metal4 ;
  RECT 3357.980 500.640 3359.100 501.760 ;
  LAYER metal3 ;
  RECT 3357.980 500.640 3359.100 501.760 ;
  LAYER metal2 ;
  RECT 3357.980 500.640 3359.100 501.760 ;
  LAYER metal1 ;
  RECT 3357.980 500.640 3359.100 501.760 ;
 END
END DIB119
PIN DOB119
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3344.960 500.640 3346.080 501.760 ;
  LAYER metal4 ;
  RECT 3344.960 500.640 3346.080 501.760 ;
  LAYER metal3 ;
  RECT 3344.960 500.640 3346.080 501.760 ;
  LAYER metal2 ;
  RECT 3344.960 500.640 3346.080 501.760 ;
  LAYER metal1 ;
  RECT 3344.960 500.640 3346.080 501.760 ;
 END
END DOB119
PIN DIB118
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3331.320 500.640 3332.440 501.760 ;
  LAYER metal4 ;
  RECT 3331.320 500.640 3332.440 501.760 ;
  LAYER metal3 ;
  RECT 3331.320 500.640 3332.440 501.760 ;
  LAYER metal2 ;
  RECT 3331.320 500.640 3332.440 501.760 ;
  LAYER metal1 ;
  RECT 3331.320 500.640 3332.440 501.760 ;
 END
END DIB118
PIN DOB118
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3317.680 500.640 3318.800 501.760 ;
  LAYER metal4 ;
  RECT 3317.680 500.640 3318.800 501.760 ;
  LAYER metal3 ;
  RECT 3317.680 500.640 3318.800 501.760 ;
  LAYER metal2 ;
  RECT 3317.680 500.640 3318.800 501.760 ;
  LAYER metal1 ;
  RECT 3317.680 500.640 3318.800 501.760 ;
 END
END DOB118
PIN DIB117
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3304.660 500.640 3305.780 501.760 ;
  LAYER metal4 ;
  RECT 3304.660 500.640 3305.780 501.760 ;
  LAYER metal3 ;
  RECT 3304.660 500.640 3305.780 501.760 ;
  LAYER metal2 ;
  RECT 3304.660 500.640 3305.780 501.760 ;
  LAYER metal1 ;
  RECT 3304.660 500.640 3305.780 501.760 ;
 END
END DIB117
PIN DOB117
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3291.020 500.640 3292.140 501.760 ;
  LAYER metal4 ;
  RECT 3291.020 500.640 3292.140 501.760 ;
  LAYER metal3 ;
  RECT 3291.020 500.640 3292.140 501.760 ;
  LAYER metal2 ;
  RECT 3291.020 500.640 3292.140 501.760 ;
  LAYER metal1 ;
  RECT 3291.020 500.640 3292.140 501.760 ;
 END
END DOB117
PIN DIB116
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3277.380 500.640 3278.500 501.760 ;
  LAYER metal4 ;
  RECT 3277.380 500.640 3278.500 501.760 ;
  LAYER metal3 ;
  RECT 3277.380 500.640 3278.500 501.760 ;
  LAYER metal2 ;
  RECT 3277.380 500.640 3278.500 501.760 ;
  LAYER metal1 ;
  RECT 3277.380 500.640 3278.500 501.760 ;
 END
END DIB116
PIN DOB116
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3264.360 500.640 3265.480 501.760 ;
  LAYER metal4 ;
  RECT 3264.360 500.640 3265.480 501.760 ;
  LAYER metal3 ;
  RECT 3264.360 500.640 3265.480 501.760 ;
  LAYER metal2 ;
  RECT 3264.360 500.640 3265.480 501.760 ;
  LAYER metal1 ;
  RECT 3264.360 500.640 3265.480 501.760 ;
 END
END DOB116
PIN DIB115
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3250.720 500.640 3251.840 501.760 ;
  LAYER metal4 ;
  RECT 3250.720 500.640 3251.840 501.760 ;
  LAYER metal3 ;
  RECT 3250.720 500.640 3251.840 501.760 ;
  LAYER metal2 ;
  RECT 3250.720 500.640 3251.840 501.760 ;
  LAYER metal1 ;
  RECT 3250.720 500.640 3251.840 501.760 ;
 END
END DIB115
PIN DOB115
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3237.080 500.640 3238.200 501.760 ;
  LAYER metal4 ;
  RECT 3237.080 500.640 3238.200 501.760 ;
  LAYER metal3 ;
  RECT 3237.080 500.640 3238.200 501.760 ;
  LAYER metal2 ;
  RECT 3237.080 500.640 3238.200 501.760 ;
  LAYER metal1 ;
  RECT 3237.080 500.640 3238.200 501.760 ;
 END
END DOB115
PIN DIB114
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3224.060 500.640 3225.180 501.760 ;
  LAYER metal4 ;
  RECT 3224.060 500.640 3225.180 501.760 ;
  LAYER metal3 ;
  RECT 3224.060 500.640 3225.180 501.760 ;
  LAYER metal2 ;
  RECT 3224.060 500.640 3225.180 501.760 ;
  LAYER metal1 ;
  RECT 3224.060 500.640 3225.180 501.760 ;
 END
END DIB114
PIN DOB114
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3210.420 500.640 3211.540 501.760 ;
  LAYER metal4 ;
  RECT 3210.420 500.640 3211.540 501.760 ;
  LAYER metal3 ;
  RECT 3210.420 500.640 3211.540 501.760 ;
  LAYER metal2 ;
  RECT 3210.420 500.640 3211.540 501.760 ;
  LAYER metal1 ;
  RECT 3210.420 500.640 3211.540 501.760 ;
 END
END DOB114
PIN DIB113
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3196.780 500.640 3197.900 501.760 ;
  LAYER metal4 ;
  RECT 3196.780 500.640 3197.900 501.760 ;
  LAYER metal3 ;
  RECT 3196.780 500.640 3197.900 501.760 ;
  LAYER metal2 ;
  RECT 3196.780 500.640 3197.900 501.760 ;
  LAYER metal1 ;
  RECT 3196.780 500.640 3197.900 501.760 ;
 END
END DIB113
PIN DOB113
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3183.760 500.640 3184.880 501.760 ;
  LAYER metal4 ;
  RECT 3183.760 500.640 3184.880 501.760 ;
  LAYER metal3 ;
  RECT 3183.760 500.640 3184.880 501.760 ;
  LAYER metal2 ;
  RECT 3183.760 500.640 3184.880 501.760 ;
  LAYER metal1 ;
  RECT 3183.760 500.640 3184.880 501.760 ;
 END
END DOB113
PIN DIB112
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3170.120 500.640 3171.240 501.760 ;
  LAYER metal4 ;
  RECT 3170.120 500.640 3171.240 501.760 ;
  LAYER metal3 ;
  RECT 3170.120 500.640 3171.240 501.760 ;
  LAYER metal2 ;
  RECT 3170.120 500.640 3171.240 501.760 ;
  LAYER metal1 ;
  RECT 3170.120 500.640 3171.240 501.760 ;
 END
END DIB112
PIN DOB112
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3156.480 500.640 3157.600 501.760 ;
  LAYER metal4 ;
  RECT 3156.480 500.640 3157.600 501.760 ;
  LAYER metal3 ;
  RECT 3156.480 500.640 3157.600 501.760 ;
  LAYER metal2 ;
  RECT 3156.480 500.640 3157.600 501.760 ;
  LAYER metal1 ;
  RECT 3156.480 500.640 3157.600 501.760 ;
 END
END DOB112
PIN DIB111
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3142.840 500.640 3143.960 501.760 ;
  LAYER metal4 ;
  RECT 3142.840 500.640 3143.960 501.760 ;
  LAYER metal3 ;
  RECT 3142.840 500.640 3143.960 501.760 ;
  LAYER metal2 ;
  RECT 3142.840 500.640 3143.960 501.760 ;
  LAYER metal1 ;
  RECT 3142.840 500.640 3143.960 501.760 ;
 END
END DIB111
PIN DOB111
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3129.820 500.640 3130.940 501.760 ;
  LAYER metal4 ;
  RECT 3129.820 500.640 3130.940 501.760 ;
  LAYER metal3 ;
  RECT 3129.820 500.640 3130.940 501.760 ;
  LAYER metal2 ;
  RECT 3129.820 500.640 3130.940 501.760 ;
  LAYER metal1 ;
  RECT 3129.820 500.640 3130.940 501.760 ;
 END
END DOB111
PIN DIB110
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3116.180 500.640 3117.300 501.760 ;
  LAYER metal4 ;
  RECT 3116.180 500.640 3117.300 501.760 ;
  LAYER metal3 ;
  RECT 3116.180 500.640 3117.300 501.760 ;
  LAYER metal2 ;
  RECT 3116.180 500.640 3117.300 501.760 ;
  LAYER metal1 ;
  RECT 3116.180 500.640 3117.300 501.760 ;
 END
END DIB110
PIN DOB110
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3102.540 500.640 3103.660 501.760 ;
  LAYER metal4 ;
  RECT 3102.540 500.640 3103.660 501.760 ;
  LAYER metal3 ;
  RECT 3102.540 500.640 3103.660 501.760 ;
  LAYER metal2 ;
  RECT 3102.540 500.640 3103.660 501.760 ;
  LAYER metal1 ;
  RECT 3102.540 500.640 3103.660 501.760 ;
 END
END DOB110
PIN DIB109
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3089.520 500.640 3090.640 501.760 ;
  LAYER metal4 ;
  RECT 3089.520 500.640 3090.640 501.760 ;
  LAYER metal3 ;
  RECT 3089.520 500.640 3090.640 501.760 ;
  LAYER metal2 ;
  RECT 3089.520 500.640 3090.640 501.760 ;
  LAYER metal1 ;
  RECT 3089.520 500.640 3090.640 501.760 ;
 END
END DIB109
PIN DOB109
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3075.880 500.640 3077.000 501.760 ;
  LAYER metal4 ;
  RECT 3075.880 500.640 3077.000 501.760 ;
  LAYER metal3 ;
  RECT 3075.880 500.640 3077.000 501.760 ;
  LAYER metal2 ;
  RECT 3075.880 500.640 3077.000 501.760 ;
  LAYER metal1 ;
  RECT 3075.880 500.640 3077.000 501.760 ;
 END
END DOB109
PIN DIB108
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3062.240 500.640 3063.360 501.760 ;
  LAYER metal4 ;
  RECT 3062.240 500.640 3063.360 501.760 ;
  LAYER metal3 ;
  RECT 3062.240 500.640 3063.360 501.760 ;
  LAYER metal2 ;
  RECT 3062.240 500.640 3063.360 501.760 ;
  LAYER metal1 ;
  RECT 3062.240 500.640 3063.360 501.760 ;
 END
END DIB108
PIN DOB108
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3049.220 500.640 3050.340 501.760 ;
  LAYER metal4 ;
  RECT 3049.220 500.640 3050.340 501.760 ;
  LAYER metal3 ;
  RECT 3049.220 500.640 3050.340 501.760 ;
  LAYER metal2 ;
  RECT 3049.220 500.640 3050.340 501.760 ;
  LAYER metal1 ;
  RECT 3049.220 500.640 3050.340 501.760 ;
 END
END DOB108
PIN DIB107
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3035.580 500.640 3036.700 501.760 ;
  LAYER metal4 ;
  RECT 3035.580 500.640 3036.700 501.760 ;
  LAYER metal3 ;
  RECT 3035.580 500.640 3036.700 501.760 ;
  LAYER metal2 ;
  RECT 3035.580 500.640 3036.700 501.760 ;
  LAYER metal1 ;
  RECT 3035.580 500.640 3036.700 501.760 ;
 END
END DIB107
PIN DOB107
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3021.940 500.640 3023.060 501.760 ;
  LAYER metal4 ;
  RECT 3021.940 500.640 3023.060 501.760 ;
  LAYER metal3 ;
  RECT 3021.940 500.640 3023.060 501.760 ;
  LAYER metal2 ;
  RECT 3021.940 500.640 3023.060 501.760 ;
  LAYER metal1 ;
  RECT 3021.940 500.640 3023.060 501.760 ;
 END
END DOB107
PIN DIB106
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3008.920 500.640 3010.040 501.760 ;
  LAYER metal4 ;
  RECT 3008.920 500.640 3010.040 501.760 ;
  LAYER metal3 ;
  RECT 3008.920 500.640 3010.040 501.760 ;
  LAYER metal2 ;
  RECT 3008.920 500.640 3010.040 501.760 ;
  LAYER metal1 ;
  RECT 3008.920 500.640 3010.040 501.760 ;
 END
END DIB106
PIN DOB106
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2995.280 500.640 2996.400 501.760 ;
  LAYER metal4 ;
  RECT 2995.280 500.640 2996.400 501.760 ;
  LAYER metal3 ;
  RECT 2995.280 500.640 2996.400 501.760 ;
  LAYER metal2 ;
  RECT 2995.280 500.640 2996.400 501.760 ;
  LAYER metal1 ;
  RECT 2995.280 500.640 2996.400 501.760 ;
 END
END DOB106
PIN DIB105
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2981.640 500.640 2982.760 501.760 ;
  LAYER metal4 ;
  RECT 2981.640 500.640 2982.760 501.760 ;
  LAYER metal3 ;
  RECT 2981.640 500.640 2982.760 501.760 ;
  LAYER metal2 ;
  RECT 2981.640 500.640 2982.760 501.760 ;
  LAYER metal1 ;
  RECT 2981.640 500.640 2982.760 501.760 ;
 END
END DIB105
PIN DOB105
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2968.620 500.640 2969.740 501.760 ;
  LAYER metal4 ;
  RECT 2968.620 500.640 2969.740 501.760 ;
  LAYER metal3 ;
  RECT 2968.620 500.640 2969.740 501.760 ;
  LAYER metal2 ;
  RECT 2968.620 500.640 2969.740 501.760 ;
  LAYER metal1 ;
  RECT 2968.620 500.640 2969.740 501.760 ;
 END
END DOB105
PIN DIB104
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2954.980 500.640 2956.100 501.760 ;
  LAYER metal4 ;
  RECT 2954.980 500.640 2956.100 501.760 ;
  LAYER metal3 ;
  RECT 2954.980 500.640 2956.100 501.760 ;
  LAYER metal2 ;
  RECT 2954.980 500.640 2956.100 501.760 ;
  LAYER metal1 ;
  RECT 2954.980 500.640 2956.100 501.760 ;
 END
END DIB104
PIN DOB104
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2941.340 500.640 2942.460 501.760 ;
  LAYER metal4 ;
  RECT 2941.340 500.640 2942.460 501.760 ;
  LAYER metal3 ;
  RECT 2941.340 500.640 2942.460 501.760 ;
  LAYER metal2 ;
  RECT 2941.340 500.640 2942.460 501.760 ;
  LAYER metal1 ;
  RECT 2941.340 500.640 2942.460 501.760 ;
 END
END DOB104
PIN DIB103
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2928.320 500.640 2929.440 501.760 ;
  LAYER metal4 ;
  RECT 2928.320 500.640 2929.440 501.760 ;
  LAYER metal3 ;
  RECT 2928.320 500.640 2929.440 501.760 ;
  LAYER metal2 ;
  RECT 2928.320 500.640 2929.440 501.760 ;
  LAYER metal1 ;
  RECT 2928.320 500.640 2929.440 501.760 ;
 END
END DIB103
PIN DOB103
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2914.680 500.640 2915.800 501.760 ;
  LAYER metal4 ;
  RECT 2914.680 500.640 2915.800 501.760 ;
  LAYER metal3 ;
  RECT 2914.680 500.640 2915.800 501.760 ;
  LAYER metal2 ;
  RECT 2914.680 500.640 2915.800 501.760 ;
  LAYER metal1 ;
  RECT 2914.680 500.640 2915.800 501.760 ;
 END
END DOB103
PIN DIB102
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2901.040 500.640 2902.160 501.760 ;
  LAYER metal4 ;
  RECT 2901.040 500.640 2902.160 501.760 ;
  LAYER metal3 ;
  RECT 2901.040 500.640 2902.160 501.760 ;
  LAYER metal2 ;
  RECT 2901.040 500.640 2902.160 501.760 ;
  LAYER metal1 ;
  RECT 2901.040 500.640 2902.160 501.760 ;
 END
END DIB102
PIN DOB102
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2888.020 500.640 2889.140 501.760 ;
  LAYER metal4 ;
  RECT 2888.020 500.640 2889.140 501.760 ;
  LAYER metal3 ;
  RECT 2888.020 500.640 2889.140 501.760 ;
  LAYER metal2 ;
  RECT 2888.020 500.640 2889.140 501.760 ;
  LAYER metal1 ;
  RECT 2888.020 500.640 2889.140 501.760 ;
 END
END DOB102
PIN DIB101
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2874.380 500.640 2875.500 501.760 ;
  LAYER metal4 ;
  RECT 2874.380 500.640 2875.500 501.760 ;
  LAYER metal3 ;
  RECT 2874.380 500.640 2875.500 501.760 ;
  LAYER metal2 ;
  RECT 2874.380 500.640 2875.500 501.760 ;
  LAYER metal1 ;
  RECT 2874.380 500.640 2875.500 501.760 ;
 END
END DIB101
PIN DOB101
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2860.740 500.640 2861.860 501.760 ;
  LAYER metal4 ;
  RECT 2860.740 500.640 2861.860 501.760 ;
  LAYER metal3 ;
  RECT 2860.740 500.640 2861.860 501.760 ;
  LAYER metal2 ;
  RECT 2860.740 500.640 2861.860 501.760 ;
  LAYER metal1 ;
  RECT 2860.740 500.640 2861.860 501.760 ;
 END
END DOB101
PIN DIB100
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2847.720 500.640 2848.840 501.760 ;
  LAYER metal4 ;
  RECT 2847.720 500.640 2848.840 501.760 ;
  LAYER metal3 ;
  RECT 2847.720 500.640 2848.840 501.760 ;
  LAYER metal2 ;
  RECT 2847.720 500.640 2848.840 501.760 ;
  LAYER metal1 ;
  RECT 2847.720 500.640 2848.840 501.760 ;
 END
END DIB100
PIN DOB100
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2834.080 500.640 2835.200 501.760 ;
  LAYER metal4 ;
  RECT 2834.080 500.640 2835.200 501.760 ;
  LAYER metal3 ;
  RECT 2834.080 500.640 2835.200 501.760 ;
  LAYER metal2 ;
  RECT 2834.080 500.640 2835.200 501.760 ;
  LAYER metal1 ;
  RECT 2834.080 500.640 2835.200 501.760 ;
 END
END DOB100
PIN DIB99
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2820.440 500.640 2821.560 501.760 ;
  LAYER metal4 ;
  RECT 2820.440 500.640 2821.560 501.760 ;
  LAYER metal3 ;
  RECT 2820.440 500.640 2821.560 501.760 ;
  LAYER metal2 ;
  RECT 2820.440 500.640 2821.560 501.760 ;
  LAYER metal1 ;
  RECT 2820.440 500.640 2821.560 501.760 ;
 END
END DIB99
PIN DOB99
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2807.420 500.640 2808.540 501.760 ;
  LAYER metal4 ;
  RECT 2807.420 500.640 2808.540 501.760 ;
  LAYER metal3 ;
  RECT 2807.420 500.640 2808.540 501.760 ;
  LAYER metal2 ;
  RECT 2807.420 500.640 2808.540 501.760 ;
  LAYER metal1 ;
  RECT 2807.420 500.640 2808.540 501.760 ;
 END
END DOB99
PIN DIB98
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2793.780 500.640 2794.900 501.760 ;
  LAYER metal4 ;
  RECT 2793.780 500.640 2794.900 501.760 ;
  LAYER metal3 ;
  RECT 2793.780 500.640 2794.900 501.760 ;
  LAYER metal2 ;
  RECT 2793.780 500.640 2794.900 501.760 ;
  LAYER metal1 ;
  RECT 2793.780 500.640 2794.900 501.760 ;
 END
END DIB98
PIN DOB98
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2780.140 500.640 2781.260 501.760 ;
  LAYER metal4 ;
  RECT 2780.140 500.640 2781.260 501.760 ;
  LAYER metal3 ;
  RECT 2780.140 500.640 2781.260 501.760 ;
  LAYER metal2 ;
  RECT 2780.140 500.640 2781.260 501.760 ;
  LAYER metal1 ;
  RECT 2780.140 500.640 2781.260 501.760 ;
 END
END DOB98
PIN DIB97
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2767.120 500.640 2768.240 501.760 ;
  LAYER metal4 ;
  RECT 2767.120 500.640 2768.240 501.760 ;
  LAYER metal3 ;
  RECT 2767.120 500.640 2768.240 501.760 ;
  LAYER metal2 ;
  RECT 2767.120 500.640 2768.240 501.760 ;
  LAYER metal1 ;
  RECT 2767.120 500.640 2768.240 501.760 ;
 END
END DIB97
PIN DOB97
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2753.480 500.640 2754.600 501.760 ;
  LAYER metal4 ;
  RECT 2753.480 500.640 2754.600 501.760 ;
  LAYER metal3 ;
  RECT 2753.480 500.640 2754.600 501.760 ;
  LAYER metal2 ;
  RECT 2753.480 500.640 2754.600 501.760 ;
  LAYER metal1 ;
  RECT 2753.480 500.640 2754.600 501.760 ;
 END
END DOB97
PIN DIB96
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2739.840 500.640 2740.960 501.760 ;
  LAYER metal4 ;
  RECT 2739.840 500.640 2740.960 501.760 ;
  LAYER metal3 ;
  RECT 2739.840 500.640 2740.960 501.760 ;
  LAYER metal2 ;
  RECT 2739.840 500.640 2740.960 501.760 ;
  LAYER metal1 ;
  RECT 2739.840 500.640 2740.960 501.760 ;
 END
END DIB96
PIN DOB96
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2726.200 500.640 2727.320 501.760 ;
  LAYER metal4 ;
  RECT 2726.200 500.640 2727.320 501.760 ;
  LAYER metal3 ;
  RECT 2726.200 500.640 2727.320 501.760 ;
  LAYER metal2 ;
  RECT 2726.200 500.640 2727.320 501.760 ;
  LAYER metal1 ;
  RECT 2726.200 500.640 2727.320 501.760 ;
 END
END DOB96
PIN DIB95
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2713.180 500.640 2714.300 501.760 ;
  LAYER metal4 ;
  RECT 2713.180 500.640 2714.300 501.760 ;
  LAYER metal3 ;
  RECT 2713.180 500.640 2714.300 501.760 ;
  LAYER metal2 ;
  RECT 2713.180 500.640 2714.300 501.760 ;
  LAYER metal1 ;
  RECT 2713.180 500.640 2714.300 501.760 ;
 END
END DIB95
PIN DOB95
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2699.540 500.640 2700.660 501.760 ;
  LAYER metal4 ;
  RECT 2699.540 500.640 2700.660 501.760 ;
  LAYER metal3 ;
  RECT 2699.540 500.640 2700.660 501.760 ;
  LAYER metal2 ;
  RECT 2699.540 500.640 2700.660 501.760 ;
  LAYER metal1 ;
  RECT 2699.540 500.640 2700.660 501.760 ;
 END
END DOB95
PIN DIB94
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2685.900 500.640 2687.020 501.760 ;
  LAYER metal4 ;
  RECT 2685.900 500.640 2687.020 501.760 ;
  LAYER metal3 ;
  RECT 2685.900 500.640 2687.020 501.760 ;
  LAYER metal2 ;
  RECT 2685.900 500.640 2687.020 501.760 ;
  LAYER metal1 ;
  RECT 2685.900 500.640 2687.020 501.760 ;
 END
END DIB94
PIN DOB94
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2672.880 500.640 2674.000 501.760 ;
  LAYER metal4 ;
  RECT 2672.880 500.640 2674.000 501.760 ;
  LAYER metal3 ;
  RECT 2672.880 500.640 2674.000 501.760 ;
  LAYER metal2 ;
  RECT 2672.880 500.640 2674.000 501.760 ;
  LAYER metal1 ;
  RECT 2672.880 500.640 2674.000 501.760 ;
 END
END DOB94
PIN DIB93
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2659.240 500.640 2660.360 501.760 ;
  LAYER metal4 ;
  RECT 2659.240 500.640 2660.360 501.760 ;
  LAYER metal3 ;
  RECT 2659.240 500.640 2660.360 501.760 ;
  LAYER metal2 ;
  RECT 2659.240 500.640 2660.360 501.760 ;
  LAYER metal1 ;
  RECT 2659.240 500.640 2660.360 501.760 ;
 END
END DIB93
PIN DOB93
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2645.600 500.640 2646.720 501.760 ;
  LAYER metal4 ;
  RECT 2645.600 500.640 2646.720 501.760 ;
  LAYER metal3 ;
  RECT 2645.600 500.640 2646.720 501.760 ;
  LAYER metal2 ;
  RECT 2645.600 500.640 2646.720 501.760 ;
  LAYER metal1 ;
  RECT 2645.600 500.640 2646.720 501.760 ;
 END
END DOB93
PIN DIB92
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2632.580 500.640 2633.700 501.760 ;
  LAYER metal4 ;
  RECT 2632.580 500.640 2633.700 501.760 ;
  LAYER metal3 ;
  RECT 2632.580 500.640 2633.700 501.760 ;
  LAYER metal2 ;
  RECT 2632.580 500.640 2633.700 501.760 ;
  LAYER metal1 ;
  RECT 2632.580 500.640 2633.700 501.760 ;
 END
END DIB92
PIN DOB92
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2618.940 500.640 2620.060 501.760 ;
  LAYER metal4 ;
  RECT 2618.940 500.640 2620.060 501.760 ;
  LAYER metal3 ;
  RECT 2618.940 500.640 2620.060 501.760 ;
  LAYER metal2 ;
  RECT 2618.940 500.640 2620.060 501.760 ;
  LAYER metal1 ;
  RECT 2618.940 500.640 2620.060 501.760 ;
 END
END DOB92
PIN DIB91
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2605.300 500.640 2606.420 501.760 ;
  LAYER metal4 ;
  RECT 2605.300 500.640 2606.420 501.760 ;
  LAYER metal3 ;
  RECT 2605.300 500.640 2606.420 501.760 ;
  LAYER metal2 ;
  RECT 2605.300 500.640 2606.420 501.760 ;
  LAYER metal1 ;
  RECT 2605.300 500.640 2606.420 501.760 ;
 END
END DIB91
PIN DOB91
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2592.280 500.640 2593.400 501.760 ;
  LAYER metal4 ;
  RECT 2592.280 500.640 2593.400 501.760 ;
  LAYER metal3 ;
  RECT 2592.280 500.640 2593.400 501.760 ;
  LAYER metal2 ;
  RECT 2592.280 500.640 2593.400 501.760 ;
  LAYER metal1 ;
  RECT 2592.280 500.640 2593.400 501.760 ;
 END
END DOB91
PIN DIB90
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2578.640 500.640 2579.760 501.760 ;
  LAYER metal4 ;
  RECT 2578.640 500.640 2579.760 501.760 ;
  LAYER metal3 ;
  RECT 2578.640 500.640 2579.760 501.760 ;
  LAYER metal2 ;
  RECT 2578.640 500.640 2579.760 501.760 ;
  LAYER metal1 ;
  RECT 2578.640 500.640 2579.760 501.760 ;
 END
END DIB90
PIN DOB90
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2565.000 500.640 2566.120 501.760 ;
  LAYER metal4 ;
  RECT 2565.000 500.640 2566.120 501.760 ;
  LAYER metal3 ;
  RECT 2565.000 500.640 2566.120 501.760 ;
  LAYER metal2 ;
  RECT 2565.000 500.640 2566.120 501.760 ;
  LAYER metal1 ;
  RECT 2565.000 500.640 2566.120 501.760 ;
 END
END DOB90
PIN DIB89
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2551.980 500.640 2553.100 501.760 ;
  LAYER metal4 ;
  RECT 2551.980 500.640 2553.100 501.760 ;
  LAYER metal3 ;
  RECT 2551.980 500.640 2553.100 501.760 ;
  LAYER metal2 ;
  RECT 2551.980 500.640 2553.100 501.760 ;
  LAYER metal1 ;
  RECT 2551.980 500.640 2553.100 501.760 ;
 END
END DIB89
PIN DOB89
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2538.340 500.640 2539.460 501.760 ;
  LAYER metal4 ;
  RECT 2538.340 500.640 2539.460 501.760 ;
  LAYER metal3 ;
  RECT 2538.340 500.640 2539.460 501.760 ;
  LAYER metal2 ;
  RECT 2538.340 500.640 2539.460 501.760 ;
  LAYER metal1 ;
  RECT 2538.340 500.640 2539.460 501.760 ;
 END
END DOB89
PIN DIB88
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2524.700 500.640 2525.820 501.760 ;
  LAYER metal4 ;
  RECT 2524.700 500.640 2525.820 501.760 ;
  LAYER metal3 ;
  RECT 2524.700 500.640 2525.820 501.760 ;
  LAYER metal2 ;
  RECT 2524.700 500.640 2525.820 501.760 ;
  LAYER metal1 ;
  RECT 2524.700 500.640 2525.820 501.760 ;
 END
END DIB88
PIN DOB88
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2511.680 500.640 2512.800 501.760 ;
  LAYER metal4 ;
  RECT 2511.680 500.640 2512.800 501.760 ;
  LAYER metal3 ;
  RECT 2511.680 500.640 2512.800 501.760 ;
  LAYER metal2 ;
  RECT 2511.680 500.640 2512.800 501.760 ;
  LAYER metal1 ;
  RECT 2511.680 500.640 2512.800 501.760 ;
 END
END DOB88
PIN DIB87
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2498.040 500.640 2499.160 501.760 ;
  LAYER metal4 ;
  RECT 2498.040 500.640 2499.160 501.760 ;
  LAYER metal3 ;
  RECT 2498.040 500.640 2499.160 501.760 ;
  LAYER metal2 ;
  RECT 2498.040 500.640 2499.160 501.760 ;
  LAYER metal1 ;
  RECT 2498.040 500.640 2499.160 501.760 ;
 END
END DIB87
PIN DOB87
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2484.400 500.640 2485.520 501.760 ;
  LAYER metal4 ;
  RECT 2484.400 500.640 2485.520 501.760 ;
  LAYER metal3 ;
  RECT 2484.400 500.640 2485.520 501.760 ;
  LAYER metal2 ;
  RECT 2484.400 500.640 2485.520 501.760 ;
  LAYER metal1 ;
  RECT 2484.400 500.640 2485.520 501.760 ;
 END
END DOB87
PIN DIB86
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2471.380 500.640 2472.500 501.760 ;
  LAYER metal4 ;
  RECT 2471.380 500.640 2472.500 501.760 ;
  LAYER metal3 ;
  RECT 2471.380 500.640 2472.500 501.760 ;
  LAYER metal2 ;
  RECT 2471.380 500.640 2472.500 501.760 ;
  LAYER metal1 ;
  RECT 2471.380 500.640 2472.500 501.760 ;
 END
END DIB86
PIN DOB86
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2457.740 500.640 2458.860 501.760 ;
  LAYER metal4 ;
  RECT 2457.740 500.640 2458.860 501.760 ;
  LAYER metal3 ;
  RECT 2457.740 500.640 2458.860 501.760 ;
  LAYER metal2 ;
  RECT 2457.740 500.640 2458.860 501.760 ;
  LAYER metal1 ;
  RECT 2457.740 500.640 2458.860 501.760 ;
 END
END DOB86
PIN DIB85
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2444.100 500.640 2445.220 501.760 ;
  LAYER metal4 ;
  RECT 2444.100 500.640 2445.220 501.760 ;
  LAYER metal3 ;
  RECT 2444.100 500.640 2445.220 501.760 ;
  LAYER metal2 ;
  RECT 2444.100 500.640 2445.220 501.760 ;
  LAYER metal1 ;
  RECT 2444.100 500.640 2445.220 501.760 ;
 END
END DIB85
PIN DOB85
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2431.080 500.640 2432.200 501.760 ;
  LAYER metal4 ;
  RECT 2431.080 500.640 2432.200 501.760 ;
  LAYER metal3 ;
  RECT 2431.080 500.640 2432.200 501.760 ;
  LAYER metal2 ;
  RECT 2431.080 500.640 2432.200 501.760 ;
  LAYER metal1 ;
  RECT 2431.080 500.640 2432.200 501.760 ;
 END
END DOB85
PIN DIB84
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2417.440 500.640 2418.560 501.760 ;
  LAYER metal4 ;
  RECT 2417.440 500.640 2418.560 501.760 ;
  LAYER metal3 ;
  RECT 2417.440 500.640 2418.560 501.760 ;
  LAYER metal2 ;
  RECT 2417.440 500.640 2418.560 501.760 ;
  LAYER metal1 ;
  RECT 2417.440 500.640 2418.560 501.760 ;
 END
END DIB84
PIN DOB84
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2403.800 500.640 2404.920 501.760 ;
  LAYER metal4 ;
  RECT 2403.800 500.640 2404.920 501.760 ;
  LAYER metal3 ;
  RECT 2403.800 500.640 2404.920 501.760 ;
  LAYER metal2 ;
  RECT 2403.800 500.640 2404.920 501.760 ;
  LAYER metal1 ;
  RECT 2403.800 500.640 2404.920 501.760 ;
 END
END DOB84
PIN DIB83
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2390.780 500.640 2391.900 501.760 ;
  LAYER metal4 ;
  RECT 2390.780 500.640 2391.900 501.760 ;
  LAYER metal3 ;
  RECT 2390.780 500.640 2391.900 501.760 ;
  LAYER metal2 ;
  RECT 2390.780 500.640 2391.900 501.760 ;
  LAYER metal1 ;
  RECT 2390.780 500.640 2391.900 501.760 ;
 END
END DIB83
PIN DOB83
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2377.140 500.640 2378.260 501.760 ;
  LAYER metal4 ;
  RECT 2377.140 500.640 2378.260 501.760 ;
  LAYER metal3 ;
  RECT 2377.140 500.640 2378.260 501.760 ;
  LAYER metal2 ;
  RECT 2377.140 500.640 2378.260 501.760 ;
  LAYER metal1 ;
  RECT 2377.140 500.640 2378.260 501.760 ;
 END
END DOB83
PIN DIB82
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2363.500 500.640 2364.620 501.760 ;
  LAYER metal4 ;
  RECT 2363.500 500.640 2364.620 501.760 ;
  LAYER metal3 ;
  RECT 2363.500 500.640 2364.620 501.760 ;
  LAYER metal2 ;
  RECT 2363.500 500.640 2364.620 501.760 ;
  LAYER metal1 ;
  RECT 2363.500 500.640 2364.620 501.760 ;
 END
END DIB82
PIN DOB82
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2350.480 500.640 2351.600 501.760 ;
  LAYER metal4 ;
  RECT 2350.480 500.640 2351.600 501.760 ;
  LAYER metal3 ;
  RECT 2350.480 500.640 2351.600 501.760 ;
  LAYER metal2 ;
  RECT 2350.480 500.640 2351.600 501.760 ;
  LAYER metal1 ;
  RECT 2350.480 500.640 2351.600 501.760 ;
 END
END DOB82
PIN DIB81
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2336.840 500.640 2337.960 501.760 ;
  LAYER metal4 ;
  RECT 2336.840 500.640 2337.960 501.760 ;
  LAYER metal3 ;
  RECT 2336.840 500.640 2337.960 501.760 ;
  LAYER metal2 ;
  RECT 2336.840 500.640 2337.960 501.760 ;
  LAYER metal1 ;
  RECT 2336.840 500.640 2337.960 501.760 ;
 END
END DIB81
PIN DOB81
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2323.200 500.640 2324.320 501.760 ;
  LAYER metal4 ;
  RECT 2323.200 500.640 2324.320 501.760 ;
  LAYER metal3 ;
  RECT 2323.200 500.640 2324.320 501.760 ;
  LAYER metal2 ;
  RECT 2323.200 500.640 2324.320 501.760 ;
  LAYER metal1 ;
  RECT 2323.200 500.640 2324.320 501.760 ;
 END
END DOB81
PIN DIB80
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2309.560 500.640 2310.680 501.760 ;
  LAYER metal4 ;
  RECT 2309.560 500.640 2310.680 501.760 ;
  LAYER metal3 ;
  RECT 2309.560 500.640 2310.680 501.760 ;
  LAYER metal2 ;
  RECT 2309.560 500.640 2310.680 501.760 ;
  LAYER metal1 ;
  RECT 2309.560 500.640 2310.680 501.760 ;
 END
END DIB80
PIN DOB80
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2296.540 500.640 2297.660 501.760 ;
  LAYER metal4 ;
  RECT 2296.540 500.640 2297.660 501.760 ;
  LAYER metal3 ;
  RECT 2296.540 500.640 2297.660 501.760 ;
  LAYER metal2 ;
  RECT 2296.540 500.640 2297.660 501.760 ;
  LAYER metal1 ;
  RECT 2296.540 500.640 2297.660 501.760 ;
 END
END DOB80
PIN DIB79
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2282.900 500.640 2284.020 501.760 ;
  LAYER metal4 ;
  RECT 2282.900 500.640 2284.020 501.760 ;
  LAYER metal3 ;
  RECT 2282.900 500.640 2284.020 501.760 ;
  LAYER metal2 ;
  RECT 2282.900 500.640 2284.020 501.760 ;
  LAYER metal1 ;
  RECT 2282.900 500.640 2284.020 501.760 ;
 END
END DIB79
PIN DOB79
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2269.260 500.640 2270.380 501.760 ;
  LAYER metal4 ;
  RECT 2269.260 500.640 2270.380 501.760 ;
  LAYER metal3 ;
  RECT 2269.260 500.640 2270.380 501.760 ;
  LAYER metal2 ;
  RECT 2269.260 500.640 2270.380 501.760 ;
  LAYER metal1 ;
  RECT 2269.260 500.640 2270.380 501.760 ;
 END
END DOB79
PIN DIB78
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2256.240 500.640 2257.360 501.760 ;
  LAYER metal4 ;
  RECT 2256.240 500.640 2257.360 501.760 ;
  LAYER metal3 ;
  RECT 2256.240 500.640 2257.360 501.760 ;
  LAYER metal2 ;
  RECT 2256.240 500.640 2257.360 501.760 ;
  LAYER metal1 ;
  RECT 2256.240 500.640 2257.360 501.760 ;
 END
END DIB78
PIN DOB78
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2242.600 500.640 2243.720 501.760 ;
  LAYER metal4 ;
  RECT 2242.600 500.640 2243.720 501.760 ;
  LAYER metal3 ;
  RECT 2242.600 500.640 2243.720 501.760 ;
  LAYER metal2 ;
  RECT 2242.600 500.640 2243.720 501.760 ;
  LAYER metal1 ;
  RECT 2242.600 500.640 2243.720 501.760 ;
 END
END DOB78
PIN DIB77
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2228.960 500.640 2230.080 501.760 ;
  LAYER metal4 ;
  RECT 2228.960 500.640 2230.080 501.760 ;
  LAYER metal3 ;
  RECT 2228.960 500.640 2230.080 501.760 ;
  LAYER metal2 ;
  RECT 2228.960 500.640 2230.080 501.760 ;
  LAYER metal1 ;
  RECT 2228.960 500.640 2230.080 501.760 ;
 END
END DIB77
PIN DOB77
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2215.940 500.640 2217.060 501.760 ;
  LAYER metal4 ;
  RECT 2215.940 500.640 2217.060 501.760 ;
  LAYER metal3 ;
  RECT 2215.940 500.640 2217.060 501.760 ;
  LAYER metal2 ;
  RECT 2215.940 500.640 2217.060 501.760 ;
  LAYER metal1 ;
  RECT 2215.940 500.640 2217.060 501.760 ;
 END
END DOB77
PIN DIB76
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2202.300 500.640 2203.420 501.760 ;
  LAYER metal4 ;
  RECT 2202.300 500.640 2203.420 501.760 ;
  LAYER metal3 ;
  RECT 2202.300 500.640 2203.420 501.760 ;
  LAYER metal2 ;
  RECT 2202.300 500.640 2203.420 501.760 ;
  LAYER metal1 ;
  RECT 2202.300 500.640 2203.420 501.760 ;
 END
END DIB76
PIN DOB76
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2188.660 500.640 2189.780 501.760 ;
  LAYER metal4 ;
  RECT 2188.660 500.640 2189.780 501.760 ;
  LAYER metal3 ;
  RECT 2188.660 500.640 2189.780 501.760 ;
  LAYER metal2 ;
  RECT 2188.660 500.640 2189.780 501.760 ;
  LAYER metal1 ;
  RECT 2188.660 500.640 2189.780 501.760 ;
 END
END DOB76
PIN DIB75
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2175.640 500.640 2176.760 501.760 ;
  LAYER metal4 ;
  RECT 2175.640 500.640 2176.760 501.760 ;
  LAYER metal3 ;
  RECT 2175.640 500.640 2176.760 501.760 ;
  LAYER metal2 ;
  RECT 2175.640 500.640 2176.760 501.760 ;
  LAYER metal1 ;
  RECT 2175.640 500.640 2176.760 501.760 ;
 END
END DIB75
PIN DOB75
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2162.000 500.640 2163.120 501.760 ;
  LAYER metal4 ;
  RECT 2162.000 500.640 2163.120 501.760 ;
  LAYER metal3 ;
  RECT 2162.000 500.640 2163.120 501.760 ;
  LAYER metal2 ;
  RECT 2162.000 500.640 2163.120 501.760 ;
  LAYER metal1 ;
  RECT 2162.000 500.640 2163.120 501.760 ;
 END
END DOB75
PIN DIB74
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2148.360 500.640 2149.480 501.760 ;
  LAYER metal4 ;
  RECT 2148.360 500.640 2149.480 501.760 ;
  LAYER metal3 ;
  RECT 2148.360 500.640 2149.480 501.760 ;
  LAYER metal2 ;
  RECT 2148.360 500.640 2149.480 501.760 ;
  LAYER metal1 ;
  RECT 2148.360 500.640 2149.480 501.760 ;
 END
END DIB74
PIN DOB74
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2135.340 500.640 2136.460 501.760 ;
  LAYER metal4 ;
  RECT 2135.340 500.640 2136.460 501.760 ;
  LAYER metal3 ;
  RECT 2135.340 500.640 2136.460 501.760 ;
  LAYER metal2 ;
  RECT 2135.340 500.640 2136.460 501.760 ;
  LAYER metal1 ;
  RECT 2135.340 500.640 2136.460 501.760 ;
 END
END DOB74
PIN DIB73
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2121.700 500.640 2122.820 501.760 ;
  LAYER metal4 ;
  RECT 2121.700 500.640 2122.820 501.760 ;
  LAYER metal3 ;
  RECT 2121.700 500.640 2122.820 501.760 ;
  LAYER metal2 ;
  RECT 2121.700 500.640 2122.820 501.760 ;
  LAYER metal1 ;
  RECT 2121.700 500.640 2122.820 501.760 ;
 END
END DIB73
PIN DOB73
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2108.060 500.640 2109.180 501.760 ;
  LAYER metal4 ;
  RECT 2108.060 500.640 2109.180 501.760 ;
  LAYER metal3 ;
  RECT 2108.060 500.640 2109.180 501.760 ;
  LAYER metal2 ;
  RECT 2108.060 500.640 2109.180 501.760 ;
  LAYER metal1 ;
  RECT 2108.060 500.640 2109.180 501.760 ;
 END
END DOB73
PIN DIB72
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2095.040 500.640 2096.160 501.760 ;
  LAYER metal4 ;
  RECT 2095.040 500.640 2096.160 501.760 ;
  LAYER metal3 ;
  RECT 2095.040 500.640 2096.160 501.760 ;
  LAYER metal2 ;
  RECT 2095.040 500.640 2096.160 501.760 ;
  LAYER metal1 ;
  RECT 2095.040 500.640 2096.160 501.760 ;
 END
END DIB72
PIN DOB72
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2081.400 500.640 2082.520 501.760 ;
  LAYER metal4 ;
  RECT 2081.400 500.640 2082.520 501.760 ;
  LAYER metal3 ;
  RECT 2081.400 500.640 2082.520 501.760 ;
  LAYER metal2 ;
  RECT 2081.400 500.640 2082.520 501.760 ;
  LAYER metal1 ;
  RECT 2081.400 500.640 2082.520 501.760 ;
 END
END DOB72
PIN DIB71
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2067.760 500.640 2068.880 501.760 ;
  LAYER metal4 ;
  RECT 2067.760 500.640 2068.880 501.760 ;
  LAYER metal3 ;
  RECT 2067.760 500.640 2068.880 501.760 ;
  LAYER metal2 ;
  RECT 2067.760 500.640 2068.880 501.760 ;
  LAYER metal1 ;
  RECT 2067.760 500.640 2068.880 501.760 ;
 END
END DIB71
PIN DOB71
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2054.740 500.640 2055.860 501.760 ;
  LAYER metal4 ;
  RECT 2054.740 500.640 2055.860 501.760 ;
  LAYER metal3 ;
  RECT 2054.740 500.640 2055.860 501.760 ;
  LAYER metal2 ;
  RECT 2054.740 500.640 2055.860 501.760 ;
  LAYER metal1 ;
  RECT 2054.740 500.640 2055.860 501.760 ;
 END
END DOB71
PIN DIB70
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2041.100 500.640 2042.220 501.760 ;
  LAYER metal4 ;
  RECT 2041.100 500.640 2042.220 501.760 ;
  LAYER metal3 ;
  RECT 2041.100 500.640 2042.220 501.760 ;
  LAYER metal2 ;
  RECT 2041.100 500.640 2042.220 501.760 ;
  LAYER metal1 ;
  RECT 2041.100 500.640 2042.220 501.760 ;
 END
END DIB70
PIN DOB70
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2027.460 500.640 2028.580 501.760 ;
  LAYER metal4 ;
  RECT 2027.460 500.640 2028.580 501.760 ;
  LAYER metal3 ;
  RECT 2027.460 500.640 2028.580 501.760 ;
  LAYER metal2 ;
  RECT 2027.460 500.640 2028.580 501.760 ;
  LAYER metal1 ;
  RECT 2027.460 500.640 2028.580 501.760 ;
 END
END DOB70
PIN DIB69
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2014.440 500.640 2015.560 501.760 ;
  LAYER metal4 ;
  RECT 2014.440 500.640 2015.560 501.760 ;
  LAYER metal3 ;
  RECT 2014.440 500.640 2015.560 501.760 ;
  LAYER metal2 ;
  RECT 2014.440 500.640 2015.560 501.760 ;
  LAYER metal1 ;
  RECT 2014.440 500.640 2015.560 501.760 ;
 END
END DIB69
PIN DOB69
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2000.800 500.640 2001.920 501.760 ;
  LAYER metal4 ;
  RECT 2000.800 500.640 2001.920 501.760 ;
  LAYER metal3 ;
  RECT 2000.800 500.640 2001.920 501.760 ;
  LAYER metal2 ;
  RECT 2000.800 500.640 2001.920 501.760 ;
  LAYER metal1 ;
  RECT 2000.800 500.640 2001.920 501.760 ;
 END
END DOB69
PIN DIB68
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1987.160 500.640 1988.280 501.760 ;
  LAYER metal4 ;
  RECT 1987.160 500.640 1988.280 501.760 ;
  LAYER metal3 ;
  RECT 1987.160 500.640 1988.280 501.760 ;
  LAYER metal2 ;
  RECT 1987.160 500.640 1988.280 501.760 ;
  LAYER metal1 ;
  RECT 1987.160 500.640 1988.280 501.760 ;
 END
END DIB68
PIN DOB68
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1974.140 500.640 1975.260 501.760 ;
  LAYER metal4 ;
  RECT 1974.140 500.640 1975.260 501.760 ;
  LAYER metal3 ;
  RECT 1974.140 500.640 1975.260 501.760 ;
  LAYER metal2 ;
  RECT 1974.140 500.640 1975.260 501.760 ;
  LAYER metal1 ;
  RECT 1974.140 500.640 1975.260 501.760 ;
 END
END DOB68
PIN DIB67
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1960.500 500.640 1961.620 501.760 ;
  LAYER metal4 ;
  RECT 1960.500 500.640 1961.620 501.760 ;
  LAYER metal3 ;
  RECT 1960.500 500.640 1961.620 501.760 ;
  LAYER metal2 ;
  RECT 1960.500 500.640 1961.620 501.760 ;
  LAYER metal1 ;
  RECT 1960.500 500.640 1961.620 501.760 ;
 END
END DIB67
PIN DOB67
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1946.860 500.640 1947.980 501.760 ;
  LAYER metal4 ;
  RECT 1946.860 500.640 1947.980 501.760 ;
  LAYER metal3 ;
  RECT 1946.860 500.640 1947.980 501.760 ;
  LAYER metal2 ;
  RECT 1946.860 500.640 1947.980 501.760 ;
  LAYER metal1 ;
  RECT 1946.860 500.640 1947.980 501.760 ;
 END
END DOB67
PIN DIB66
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1933.840 500.640 1934.960 501.760 ;
  LAYER metal4 ;
  RECT 1933.840 500.640 1934.960 501.760 ;
  LAYER metal3 ;
  RECT 1933.840 500.640 1934.960 501.760 ;
  LAYER metal2 ;
  RECT 1933.840 500.640 1934.960 501.760 ;
  LAYER metal1 ;
  RECT 1933.840 500.640 1934.960 501.760 ;
 END
END DIB66
PIN DOB66
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1920.200 500.640 1921.320 501.760 ;
  LAYER metal4 ;
  RECT 1920.200 500.640 1921.320 501.760 ;
  LAYER metal3 ;
  RECT 1920.200 500.640 1921.320 501.760 ;
  LAYER metal2 ;
  RECT 1920.200 500.640 1921.320 501.760 ;
  LAYER metal1 ;
  RECT 1920.200 500.640 1921.320 501.760 ;
 END
END DOB66
PIN DIB65
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1906.560 500.640 1907.680 501.760 ;
  LAYER metal4 ;
  RECT 1906.560 500.640 1907.680 501.760 ;
  LAYER metal3 ;
  RECT 1906.560 500.640 1907.680 501.760 ;
  LAYER metal2 ;
  RECT 1906.560 500.640 1907.680 501.760 ;
  LAYER metal1 ;
  RECT 1906.560 500.640 1907.680 501.760 ;
 END
END DIB65
PIN DOB65
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1892.920 500.640 1894.040 501.760 ;
  LAYER metal4 ;
  RECT 1892.920 500.640 1894.040 501.760 ;
  LAYER metal3 ;
  RECT 1892.920 500.640 1894.040 501.760 ;
  LAYER metal2 ;
  RECT 1892.920 500.640 1894.040 501.760 ;
  LAYER metal1 ;
  RECT 1892.920 500.640 1894.040 501.760 ;
 END
END DOB65
PIN DIB64
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1879.900 500.640 1881.020 501.760 ;
  LAYER metal4 ;
  RECT 1879.900 500.640 1881.020 501.760 ;
  LAYER metal3 ;
  RECT 1879.900 500.640 1881.020 501.760 ;
  LAYER metal2 ;
  RECT 1879.900 500.640 1881.020 501.760 ;
  LAYER metal1 ;
  RECT 1879.900 500.640 1881.020 501.760 ;
 END
END DIB64
PIN DOB64
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1866.260 500.640 1867.380 501.760 ;
  LAYER metal4 ;
  RECT 1866.260 500.640 1867.380 501.760 ;
  LAYER metal3 ;
  RECT 1866.260 500.640 1867.380 501.760 ;
  LAYER metal2 ;
  RECT 1866.260 500.640 1867.380 501.760 ;
  LAYER metal1 ;
  RECT 1866.260 500.640 1867.380 501.760 ;
 END
END DOB64
PIN OEB
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1839.600 500.640 1840.720 501.760 ;
  LAYER metal4 ;
  RECT 1839.600 500.640 1840.720 501.760 ;
  LAYER metal3 ;
  RECT 1839.600 500.640 1840.720 501.760 ;
  LAYER metal2 ;
  RECT 1839.600 500.640 1840.720 501.760 ;
  LAYER metal1 ;
  RECT 1839.600 500.640 1840.720 501.760 ;
 END
END OEB
PIN CKB
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1826.580 500.640 1827.700 501.760 ;
  LAYER metal4 ;
  RECT 1826.580 500.640 1827.700 501.760 ;
  LAYER metal3 ;
  RECT 1826.580 500.640 1827.700 501.760 ;
  LAYER metal2 ;
  RECT 1826.580 500.640 1827.700 501.760 ;
  LAYER metal1 ;
  RECT 1826.580 500.640 1827.700 501.760 ;
 END
END CKB
PIN CSB
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1824.720 500.640 1825.840 501.760 ;
  LAYER metal4 ;
  RECT 1824.720 500.640 1825.840 501.760 ;
  LAYER metal3 ;
  RECT 1824.720 500.640 1825.840 501.760 ;
  LAYER metal2 ;
  RECT 1824.720 500.640 1825.840 501.760 ;
  LAYER metal1 ;
  RECT 1824.720 500.640 1825.840 501.760 ;
 END
END CSB
PIN WEBN
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1821.620 500.640 1822.740 501.760 ;
  LAYER metal4 ;
  RECT 1821.620 500.640 1822.740 501.760 ;
  LAYER metal3 ;
  RECT 1821.620 500.640 1822.740 501.760 ;
  LAYER metal2 ;
  RECT 1821.620 500.640 1822.740 501.760 ;
  LAYER metal1 ;
  RECT 1821.620 500.640 1822.740 501.760 ;
 END
END WEBN
PIN B2
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1817.900 500.640 1819.020 501.760 ;
  LAYER metal4 ;
  RECT 1817.900 500.640 1819.020 501.760 ;
  LAYER metal3 ;
  RECT 1817.900 500.640 1819.020 501.760 ;
  LAYER metal2 ;
  RECT 1817.900 500.640 1819.020 501.760 ;
  LAYER metal1 ;
  RECT 1817.900 500.640 1819.020 501.760 ;
 END
END B2
PIN B1
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1812.940 500.640 1814.060 501.760 ;
  LAYER metal4 ;
  RECT 1812.940 500.640 1814.060 501.760 ;
  LAYER metal3 ;
  RECT 1812.940 500.640 1814.060 501.760 ;
  LAYER metal2 ;
  RECT 1812.940 500.640 1814.060 501.760 ;
  LAYER metal1 ;
  RECT 1812.940 500.640 1814.060 501.760 ;
 END
END B1
PIN B0
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1810.460 500.640 1811.580 501.760 ;
  LAYER metal4 ;
  RECT 1810.460 500.640 1811.580 501.760 ;
  LAYER metal3 ;
  RECT 1810.460 500.640 1811.580 501.760 ;
  LAYER metal2 ;
  RECT 1810.460 500.640 1811.580 501.760 ;
  LAYER metal1 ;
  RECT 1810.460 500.640 1811.580 501.760 ;
 END
END B0
PIN B5
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1801.780 500.640 1802.900 501.760 ;
  LAYER metal4 ;
  RECT 1801.780 500.640 1802.900 501.760 ;
  LAYER metal3 ;
  RECT 1801.780 500.640 1802.900 501.760 ;
  LAYER metal2 ;
  RECT 1801.780 500.640 1802.900 501.760 ;
  LAYER metal1 ;
  RECT 1801.780 500.640 1802.900 501.760 ;
 END
END B5
PIN B4
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1796.200 500.640 1797.320 501.760 ;
  LAYER metal4 ;
  RECT 1796.200 500.640 1797.320 501.760 ;
  LAYER metal3 ;
  RECT 1796.200 500.640 1797.320 501.760 ;
  LAYER metal2 ;
  RECT 1796.200 500.640 1797.320 501.760 ;
  LAYER metal1 ;
  RECT 1796.200 500.640 1797.320 501.760 ;
 END
END B4
PIN B3
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1790.620 500.640 1791.740 501.760 ;
  LAYER metal4 ;
  RECT 1790.620 500.640 1791.740 501.760 ;
  LAYER metal3 ;
  RECT 1790.620 500.640 1791.740 501.760 ;
  LAYER metal2 ;
  RECT 1790.620 500.640 1791.740 501.760 ;
  LAYER metal1 ;
  RECT 1790.620 500.640 1791.740 501.760 ;
 END
END B3
PIN B8
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1777.600 500.640 1778.720 501.760 ;
  LAYER metal4 ;
  RECT 1777.600 500.640 1778.720 501.760 ;
  LAYER metal3 ;
  RECT 1777.600 500.640 1778.720 501.760 ;
  LAYER metal2 ;
  RECT 1777.600 500.640 1778.720 501.760 ;
  LAYER metal1 ;
  RECT 1777.600 500.640 1778.720 501.760 ;
 END
END B8
PIN B7
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1772.020 500.640 1773.140 501.760 ;
  LAYER metal4 ;
  RECT 1772.020 500.640 1773.140 501.760 ;
  LAYER metal3 ;
  RECT 1772.020 500.640 1773.140 501.760 ;
  LAYER metal2 ;
  RECT 1772.020 500.640 1773.140 501.760 ;
  LAYER metal1 ;
  RECT 1772.020 500.640 1773.140 501.760 ;
 END
END B7
PIN B6
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1766.440 500.640 1767.560 501.760 ;
  LAYER metal4 ;
  RECT 1766.440 500.640 1767.560 501.760 ;
  LAYER metal3 ;
  RECT 1766.440 500.640 1767.560 501.760 ;
  LAYER metal2 ;
  RECT 1766.440 500.640 1767.560 501.760 ;
  LAYER metal1 ;
  RECT 1766.440 500.640 1767.560 501.760 ;
 END
END B6
PIN B9
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1741.640 500.640 1742.760 501.760 ;
  LAYER metal4 ;
  RECT 1741.640 500.640 1742.760 501.760 ;
  LAYER metal3 ;
  RECT 1741.640 500.640 1742.760 501.760 ;
  LAYER metal2 ;
  RECT 1741.640 500.640 1742.760 501.760 ;
  LAYER metal1 ;
  RECT 1741.640 500.640 1742.760 501.760 ;
 END
END B9
PIN DIB63
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1719.320 500.640 1720.440 501.760 ;
  LAYER metal4 ;
  RECT 1719.320 500.640 1720.440 501.760 ;
  LAYER metal3 ;
  RECT 1719.320 500.640 1720.440 501.760 ;
  LAYER metal2 ;
  RECT 1719.320 500.640 1720.440 501.760 ;
  LAYER metal1 ;
  RECT 1719.320 500.640 1720.440 501.760 ;
 END
END DIB63
PIN DOB63
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1706.300 500.640 1707.420 501.760 ;
  LAYER metal4 ;
  RECT 1706.300 500.640 1707.420 501.760 ;
  LAYER metal3 ;
  RECT 1706.300 500.640 1707.420 501.760 ;
  LAYER metal2 ;
  RECT 1706.300 500.640 1707.420 501.760 ;
  LAYER metal1 ;
  RECT 1706.300 500.640 1707.420 501.760 ;
 END
END DOB63
PIN DIB62
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1692.660 500.640 1693.780 501.760 ;
  LAYER metal4 ;
  RECT 1692.660 500.640 1693.780 501.760 ;
  LAYER metal3 ;
  RECT 1692.660 500.640 1693.780 501.760 ;
  LAYER metal2 ;
  RECT 1692.660 500.640 1693.780 501.760 ;
  LAYER metal1 ;
  RECT 1692.660 500.640 1693.780 501.760 ;
 END
END DIB62
PIN DOB62
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1679.020 500.640 1680.140 501.760 ;
  LAYER metal4 ;
  RECT 1679.020 500.640 1680.140 501.760 ;
  LAYER metal3 ;
  RECT 1679.020 500.640 1680.140 501.760 ;
  LAYER metal2 ;
  RECT 1679.020 500.640 1680.140 501.760 ;
  LAYER metal1 ;
  RECT 1679.020 500.640 1680.140 501.760 ;
 END
END DOB62
PIN DIB61
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1666.000 500.640 1667.120 501.760 ;
  LAYER metal4 ;
  RECT 1666.000 500.640 1667.120 501.760 ;
  LAYER metal3 ;
  RECT 1666.000 500.640 1667.120 501.760 ;
  LAYER metal2 ;
  RECT 1666.000 500.640 1667.120 501.760 ;
  LAYER metal1 ;
  RECT 1666.000 500.640 1667.120 501.760 ;
 END
END DIB61
PIN DOB61
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1652.360 500.640 1653.480 501.760 ;
  LAYER metal4 ;
  RECT 1652.360 500.640 1653.480 501.760 ;
  LAYER metal3 ;
  RECT 1652.360 500.640 1653.480 501.760 ;
  LAYER metal2 ;
  RECT 1652.360 500.640 1653.480 501.760 ;
  LAYER metal1 ;
  RECT 1652.360 500.640 1653.480 501.760 ;
 END
END DOB61
PIN DIB60
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1638.720 500.640 1639.840 501.760 ;
  LAYER metal4 ;
  RECT 1638.720 500.640 1639.840 501.760 ;
  LAYER metal3 ;
  RECT 1638.720 500.640 1639.840 501.760 ;
  LAYER metal2 ;
  RECT 1638.720 500.640 1639.840 501.760 ;
  LAYER metal1 ;
  RECT 1638.720 500.640 1639.840 501.760 ;
 END
END DIB60
PIN DOB60
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1625.700 500.640 1626.820 501.760 ;
  LAYER metal4 ;
  RECT 1625.700 500.640 1626.820 501.760 ;
  LAYER metal3 ;
  RECT 1625.700 500.640 1626.820 501.760 ;
  LAYER metal2 ;
  RECT 1625.700 500.640 1626.820 501.760 ;
  LAYER metal1 ;
  RECT 1625.700 500.640 1626.820 501.760 ;
 END
END DOB60
PIN DIB59
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1612.060 500.640 1613.180 501.760 ;
  LAYER metal4 ;
  RECT 1612.060 500.640 1613.180 501.760 ;
  LAYER metal3 ;
  RECT 1612.060 500.640 1613.180 501.760 ;
  LAYER metal2 ;
  RECT 1612.060 500.640 1613.180 501.760 ;
  LAYER metal1 ;
  RECT 1612.060 500.640 1613.180 501.760 ;
 END
END DIB59
PIN DOB59
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1598.420 500.640 1599.540 501.760 ;
  LAYER metal4 ;
  RECT 1598.420 500.640 1599.540 501.760 ;
  LAYER metal3 ;
  RECT 1598.420 500.640 1599.540 501.760 ;
  LAYER metal2 ;
  RECT 1598.420 500.640 1599.540 501.760 ;
  LAYER metal1 ;
  RECT 1598.420 500.640 1599.540 501.760 ;
 END
END DOB59
PIN DIB58
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1585.400 500.640 1586.520 501.760 ;
  LAYER metal4 ;
  RECT 1585.400 500.640 1586.520 501.760 ;
  LAYER metal3 ;
  RECT 1585.400 500.640 1586.520 501.760 ;
  LAYER metal2 ;
  RECT 1585.400 500.640 1586.520 501.760 ;
  LAYER metal1 ;
  RECT 1585.400 500.640 1586.520 501.760 ;
 END
END DIB58
PIN DOB58
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1571.760 500.640 1572.880 501.760 ;
  LAYER metal4 ;
  RECT 1571.760 500.640 1572.880 501.760 ;
  LAYER metal3 ;
  RECT 1571.760 500.640 1572.880 501.760 ;
  LAYER metal2 ;
  RECT 1571.760 500.640 1572.880 501.760 ;
  LAYER metal1 ;
  RECT 1571.760 500.640 1572.880 501.760 ;
 END
END DOB58
PIN DIB57
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1558.120 500.640 1559.240 501.760 ;
  LAYER metal4 ;
  RECT 1558.120 500.640 1559.240 501.760 ;
  LAYER metal3 ;
  RECT 1558.120 500.640 1559.240 501.760 ;
  LAYER metal2 ;
  RECT 1558.120 500.640 1559.240 501.760 ;
  LAYER metal1 ;
  RECT 1558.120 500.640 1559.240 501.760 ;
 END
END DIB57
PIN DOB57
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1545.100 500.640 1546.220 501.760 ;
  LAYER metal4 ;
  RECT 1545.100 500.640 1546.220 501.760 ;
  LAYER metal3 ;
  RECT 1545.100 500.640 1546.220 501.760 ;
  LAYER metal2 ;
  RECT 1545.100 500.640 1546.220 501.760 ;
  LAYER metal1 ;
  RECT 1545.100 500.640 1546.220 501.760 ;
 END
END DOB57
PIN DIB56
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1531.460 500.640 1532.580 501.760 ;
  LAYER metal4 ;
  RECT 1531.460 500.640 1532.580 501.760 ;
  LAYER metal3 ;
  RECT 1531.460 500.640 1532.580 501.760 ;
  LAYER metal2 ;
  RECT 1531.460 500.640 1532.580 501.760 ;
  LAYER metal1 ;
  RECT 1531.460 500.640 1532.580 501.760 ;
 END
END DIB56
PIN DOB56
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1517.820 500.640 1518.940 501.760 ;
  LAYER metal4 ;
  RECT 1517.820 500.640 1518.940 501.760 ;
  LAYER metal3 ;
  RECT 1517.820 500.640 1518.940 501.760 ;
  LAYER metal2 ;
  RECT 1517.820 500.640 1518.940 501.760 ;
  LAYER metal1 ;
  RECT 1517.820 500.640 1518.940 501.760 ;
 END
END DOB56
PIN DIB55
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1504.800 500.640 1505.920 501.760 ;
  LAYER metal4 ;
  RECT 1504.800 500.640 1505.920 501.760 ;
  LAYER metal3 ;
  RECT 1504.800 500.640 1505.920 501.760 ;
  LAYER metal2 ;
  RECT 1504.800 500.640 1505.920 501.760 ;
  LAYER metal1 ;
  RECT 1504.800 500.640 1505.920 501.760 ;
 END
END DIB55
PIN DOB55
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1491.160 500.640 1492.280 501.760 ;
  LAYER metal4 ;
  RECT 1491.160 500.640 1492.280 501.760 ;
  LAYER metal3 ;
  RECT 1491.160 500.640 1492.280 501.760 ;
  LAYER metal2 ;
  RECT 1491.160 500.640 1492.280 501.760 ;
  LAYER metal1 ;
  RECT 1491.160 500.640 1492.280 501.760 ;
 END
END DOB55
PIN DIB54
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1477.520 500.640 1478.640 501.760 ;
  LAYER metal4 ;
  RECT 1477.520 500.640 1478.640 501.760 ;
  LAYER metal3 ;
  RECT 1477.520 500.640 1478.640 501.760 ;
  LAYER metal2 ;
  RECT 1477.520 500.640 1478.640 501.760 ;
  LAYER metal1 ;
  RECT 1477.520 500.640 1478.640 501.760 ;
 END
END DIB54
PIN DOB54
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1464.500 500.640 1465.620 501.760 ;
  LAYER metal4 ;
  RECT 1464.500 500.640 1465.620 501.760 ;
  LAYER metal3 ;
  RECT 1464.500 500.640 1465.620 501.760 ;
  LAYER metal2 ;
  RECT 1464.500 500.640 1465.620 501.760 ;
  LAYER metal1 ;
  RECT 1464.500 500.640 1465.620 501.760 ;
 END
END DOB54
PIN DIB53
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1450.860 500.640 1451.980 501.760 ;
  LAYER metal4 ;
  RECT 1450.860 500.640 1451.980 501.760 ;
  LAYER metal3 ;
  RECT 1450.860 500.640 1451.980 501.760 ;
  LAYER metal2 ;
  RECT 1450.860 500.640 1451.980 501.760 ;
  LAYER metal1 ;
  RECT 1450.860 500.640 1451.980 501.760 ;
 END
END DIB53
PIN DOB53
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1437.220 500.640 1438.340 501.760 ;
  LAYER metal4 ;
  RECT 1437.220 500.640 1438.340 501.760 ;
  LAYER metal3 ;
  RECT 1437.220 500.640 1438.340 501.760 ;
  LAYER metal2 ;
  RECT 1437.220 500.640 1438.340 501.760 ;
  LAYER metal1 ;
  RECT 1437.220 500.640 1438.340 501.760 ;
 END
END DOB53
PIN DIB52
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1424.200 500.640 1425.320 501.760 ;
  LAYER metal4 ;
  RECT 1424.200 500.640 1425.320 501.760 ;
  LAYER metal3 ;
  RECT 1424.200 500.640 1425.320 501.760 ;
  LAYER metal2 ;
  RECT 1424.200 500.640 1425.320 501.760 ;
  LAYER metal1 ;
  RECT 1424.200 500.640 1425.320 501.760 ;
 END
END DIB52
PIN DOB52
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1410.560 500.640 1411.680 501.760 ;
  LAYER metal4 ;
  RECT 1410.560 500.640 1411.680 501.760 ;
  LAYER metal3 ;
  RECT 1410.560 500.640 1411.680 501.760 ;
  LAYER metal2 ;
  RECT 1410.560 500.640 1411.680 501.760 ;
  LAYER metal1 ;
  RECT 1410.560 500.640 1411.680 501.760 ;
 END
END DOB52
PIN DIB51
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1396.920 500.640 1398.040 501.760 ;
  LAYER metal4 ;
  RECT 1396.920 500.640 1398.040 501.760 ;
  LAYER metal3 ;
  RECT 1396.920 500.640 1398.040 501.760 ;
  LAYER metal2 ;
  RECT 1396.920 500.640 1398.040 501.760 ;
  LAYER metal1 ;
  RECT 1396.920 500.640 1398.040 501.760 ;
 END
END DIB51
PIN DOB51
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1383.900 500.640 1385.020 501.760 ;
  LAYER metal4 ;
  RECT 1383.900 500.640 1385.020 501.760 ;
  LAYER metal3 ;
  RECT 1383.900 500.640 1385.020 501.760 ;
  LAYER metal2 ;
  RECT 1383.900 500.640 1385.020 501.760 ;
  LAYER metal1 ;
  RECT 1383.900 500.640 1385.020 501.760 ;
 END
END DOB51
PIN DIB50
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1370.260 500.640 1371.380 501.760 ;
  LAYER metal4 ;
  RECT 1370.260 500.640 1371.380 501.760 ;
  LAYER metal3 ;
  RECT 1370.260 500.640 1371.380 501.760 ;
  LAYER metal2 ;
  RECT 1370.260 500.640 1371.380 501.760 ;
  LAYER metal1 ;
  RECT 1370.260 500.640 1371.380 501.760 ;
 END
END DIB50
PIN DOB50
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1356.620 500.640 1357.740 501.760 ;
  LAYER metal4 ;
  RECT 1356.620 500.640 1357.740 501.760 ;
  LAYER metal3 ;
  RECT 1356.620 500.640 1357.740 501.760 ;
  LAYER metal2 ;
  RECT 1356.620 500.640 1357.740 501.760 ;
  LAYER metal1 ;
  RECT 1356.620 500.640 1357.740 501.760 ;
 END
END DOB50
PIN DIB49
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1343.600 500.640 1344.720 501.760 ;
  LAYER metal4 ;
  RECT 1343.600 500.640 1344.720 501.760 ;
  LAYER metal3 ;
  RECT 1343.600 500.640 1344.720 501.760 ;
  LAYER metal2 ;
  RECT 1343.600 500.640 1344.720 501.760 ;
  LAYER metal1 ;
  RECT 1343.600 500.640 1344.720 501.760 ;
 END
END DIB49
PIN DOB49
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1329.960 500.640 1331.080 501.760 ;
  LAYER metal4 ;
  RECT 1329.960 500.640 1331.080 501.760 ;
  LAYER metal3 ;
  RECT 1329.960 500.640 1331.080 501.760 ;
  LAYER metal2 ;
  RECT 1329.960 500.640 1331.080 501.760 ;
  LAYER metal1 ;
  RECT 1329.960 500.640 1331.080 501.760 ;
 END
END DOB49
PIN DIB48
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1316.320 500.640 1317.440 501.760 ;
  LAYER metal4 ;
  RECT 1316.320 500.640 1317.440 501.760 ;
  LAYER metal3 ;
  RECT 1316.320 500.640 1317.440 501.760 ;
  LAYER metal2 ;
  RECT 1316.320 500.640 1317.440 501.760 ;
  LAYER metal1 ;
  RECT 1316.320 500.640 1317.440 501.760 ;
 END
END DIB48
PIN DOB48
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1302.680 500.640 1303.800 501.760 ;
  LAYER metal4 ;
  RECT 1302.680 500.640 1303.800 501.760 ;
  LAYER metal3 ;
  RECT 1302.680 500.640 1303.800 501.760 ;
  LAYER metal2 ;
  RECT 1302.680 500.640 1303.800 501.760 ;
  LAYER metal1 ;
  RECT 1302.680 500.640 1303.800 501.760 ;
 END
END DOB48
PIN DIB47
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1289.660 500.640 1290.780 501.760 ;
  LAYER metal4 ;
  RECT 1289.660 500.640 1290.780 501.760 ;
  LAYER metal3 ;
  RECT 1289.660 500.640 1290.780 501.760 ;
  LAYER metal2 ;
  RECT 1289.660 500.640 1290.780 501.760 ;
  LAYER metal1 ;
  RECT 1289.660 500.640 1290.780 501.760 ;
 END
END DIB47
PIN DOB47
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1276.020 500.640 1277.140 501.760 ;
  LAYER metal4 ;
  RECT 1276.020 500.640 1277.140 501.760 ;
  LAYER metal3 ;
  RECT 1276.020 500.640 1277.140 501.760 ;
  LAYER metal2 ;
  RECT 1276.020 500.640 1277.140 501.760 ;
  LAYER metal1 ;
  RECT 1276.020 500.640 1277.140 501.760 ;
 END
END DOB47
PIN DIB46
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1262.380 500.640 1263.500 501.760 ;
  LAYER metal4 ;
  RECT 1262.380 500.640 1263.500 501.760 ;
  LAYER metal3 ;
  RECT 1262.380 500.640 1263.500 501.760 ;
  LAYER metal2 ;
  RECT 1262.380 500.640 1263.500 501.760 ;
  LAYER metal1 ;
  RECT 1262.380 500.640 1263.500 501.760 ;
 END
END DIB46
PIN DOB46
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1249.360 500.640 1250.480 501.760 ;
  LAYER metal4 ;
  RECT 1249.360 500.640 1250.480 501.760 ;
  LAYER metal3 ;
  RECT 1249.360 500.640 1250.480 501.760 ;
  LAYER metal2 ;
  RECT 1249.360 500.640 1250.480 501.760 ;
  LAYER metal1 ;
  RECT 1249.360 500.640 1250.480 501.760 ;
 END
END DOB46
PIN DIB45
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1235.720 500.640 1236.840 501.760 ;
  LAYER metal4 ;
  RECT 1235.720 500.640 1236.840 501.760 ;
  LAYER metal3 ;
  RECT 1235.720 500.640 1236.840 501.760 ;
  LAYER metal2 ;
  RECT 1235.720 500.640 1236.840 501.760 ;
  LAYER metal1 ;
  RECT 1235.720 500.640 1236.840 501.760 ;
 END
END DIB45
PIN DOB45
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1222.080 500.640 1223.200 501.760 ;
  LAYER metal4 ;
  RECT 1222.080 500.640 1223.200 501.760 ;
  LAYER metal3 ;
  RECT 1222.080 500.640 1223.200 501.760 ;
  LAYER metal2 ;
  RECT 1222.080 500.640 1223.200 501.760 ;
  LAYER metal1 ;
  RECT 1222.080 500.640 1223.200 501.760 ;
 END
END DOB45
PIN DIB44
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1209.060 500.640 1210.180 501.760 ;
  LAYER metal4 ;
  RECT 1209.060 500.640 1210.180 501.760 ;
  LAYER metal3 ;
  RECT 1209.060 500.640 1210.180 501.760 ;
  LAYER metal2 ;
  RECT 1209.060 500.640 1210.180 501.760 ;
  LAYER metal1 ;
  RECT 1209.060 500.640 1210.180 501.760 ;
 END
END DIB44
PIN DOB44
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1195.420 500.640 1196.540 501.760 ;
  LAYER metal4 ;
  RECT 1195.420 500.640 1196.540 501.760 ;
  LAYER metal3 ;
  RECT 1195.420 500.640 1196.540 501.760 ;
  LAYER metal2 ;
  RECT 1195.420 500.640 1196.540 501.760 ;
  LAYER metal1 ;
  RECT 1195.420 500.640 1196.540 501.760 ;
 END
END DOB44
PIN DIB43
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1181.780 500.640 1182.900 501.760 ;
  LAYER metal4 ;
  RECT 1181.780 500.640 1182.900 501.760 ;
  LAYER metal3 ;
  RECT 1181.780 500.640 1182.900 501.760 ;
  LAYER metal2 ;
  RECT 1181.780 500.640 1182.900 501.760 ;
  LAYER metal1 ;
  RECT 1181.780 500.640 1182.900 501.760 ;
 END
END DIB43
PIN DOB43
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1168.760 500.640 1169.880 501.760 ;
  LAYER metal4 ;
  RECT 1168.760 500.640 1169.880 501.760 ;
  LAYER metal3 ;
  RECT 1168.760 500.640 1169.880 501.760 ;
  LAYER metal2 ;
  RECT 1168.760 500.640 1169.880 501.760 ;
  LAYER metal1 ;
  RECT 1168.760 500.640 1169.880 501.760 ;
 END
END DOB43
PIN DIB42
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1155.120 500.640 1156.240 501.760 ;
  LAYER metal4 ;
  RECT 1155.120 500.640 1156.240 501.760 ;
  LAYER metal3 ;
  RECT 1155.120 500.640 1156.240 501.760 ;
  LAYER metal2 ;
  RECT 1155.120 500.640 1156.240 501.760 ;
  LAYER metal1 ;
  RECT 1155.120 500.640 1156.240 501.760 ;
 END
END DIB42
PIN DOB42
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1141.480 500.640 1142.600 501.760 ;
  LAYER metal4 ;
  RECT 1141.480 500.640 1142.600 501.760 ;
  LAYER metal3 ;
  RECT 1141.480 500.640 1142.600 501.760 ;
  LAYER metal2 ;
  RECT 1141.480 500.640 1142.600 501.760 ;
  LAYER metal1 ;
  RECT 1141.480 500.640 1142.600 501.760 ;
 END
END DOB42
PIN DIB41
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1128.460 500.640 1129.580 501.760 ;
  LAYER metal4 ;
  RECT 1128.460 500.640 1129.580 501.760 ;
  LAYER metal3 ;
  RECT 1128.460 500.640 1129.580 501.760 ;
  LAYER metal2 ;
  RECT 1128.460 500.640 1129.580 501.760 ;
  LAYER metal1 ;
  RECT 1128.460 500.640 1129.580 501.760 ;
 END
END DIB41
PIN DOB41
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1114.820 500.640 1115.940 501.760 ;
  LAYER metal4 ;
  RECT 1114.820 500.640 1115.940 501.760 ;
  LAYER metal3 ;
  RECT 1114.820 500.640 1115.940 501.760 ;
  LAYER metal2 ;
  RECT 1114.820 500.640 1115.940 501.760 ;
  LAYER metal1 ;
  RECT 1114.820 500.640 1115.940 501.760 ;
 END
END DOB41
PIN DIB40
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1101.180 500.640 1102.300 501.760 ;
  LAYER metal4 ;
  RECT 1101.180 500.640 1102.300 501.760 ;
  LAYER metal3 ;
  RECT 1101.180 500.640 1102.300 501.760 ;
  LAYER metal2 ;
  RECT 1101.180 500.640 1102.300 501.760 ;
  LAYER metal1 ;
  RECT 1101.180 500.640 1102.300 501.760 ;
 END
END DIB40
PIN DOB40
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1088.160 500.640 1089.280 501.760 ;
  LAYER metal4 ;
  RECT 1088.160 500.640 1089.280 501.760 ;
  LAYER metal3 ;
  RECT 1088.160 500.640 1089.280 501.760 ;
  LAYER metal2 ;
  RECT 1088.160 500.640 1089.280 501.760 ;
  LAYER metal1 ;
  RECT 1088.160 500.640 1089.280 501.760 ;
 END
END DOB40
PIN DIB39
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1074.520 500.640 1075.640 501.760 ;
  LAYER metal4 ;
  RECT 1074.520 500.640 1075.640 501.760 ;
  LAYER metal3 ;
  RECT 1074.520 500.640 1075.640 501.760 ;
  LAYER metal2 ;
  RECT 1074.520 500.640 1075.640 501.760 ;
  LAYER metal1 ;
  RECT 1074.520 500.640 1075.640 501.760 ;
 END
END DIB39
PIN DOB39
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1060.880 500.640 1062.000 501.760 ;
  LAYER metal4 ;
  RECT 1060.880 500.640 1062.000 501.760 ;
  LAYER metal3 ;
  RECT 1060.880 500.640 1062.000 501.760 ;
  LAYER metal2 ;
  RECT 1060.880 500.640 1062.000 501.760 ;
  LAYER metal1 ;
  RECT 1060.880 500.640 1062.000 501.760 ;
 END
END DOB39
PIN DIB38
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1047.860 500.640 1048.980 501.760 ;
  LAYER metal4 ;
  RECT 1047.860 500.640 1048.980 501.760 ;
  LAYER metal3 ;
  RECT 1047.860 500.640 1048.980 501.760 ;
  LAYER metal2 ;
  RECT 1047.860 500.640 1048.980 501.760 ;
  LAYER metal1 ;
  RECT 1047.860 500.640 1048.980 501.760 ;
 END
END DIB38
PIN DOB38
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1034.220 500.640 1035.340 501.760 ;
  LAYER metal4 ;
  RECT 1034.220 500.640 1035.340 501.760 ;
  LAYER metal3 ;
  RECT 1034.220 500.640 1035.340 501.760 ;
  LAYER metal2 ;
  RECT 1034.220 500.640 1035.340 501.760 ;
  LAYER metal1 ;
  RECT 1034.220 500.640 1035.340 501.760 ;
 END
END DOB38
PIN DIB37
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1020.580 500.640 1021.700 501.760 ;
  LAYER metal4 ;
  RECT 1020.580 500.640 1021.700 501.760 ;
  LAYER metal3 ;
  RECT 1020.580 500.640 1021.700 501.760 ;
  LAYER metal2 ;
  RECT 1020.580 500.640 1021.700 501.760 ;
  LAYER metal1 ;
  RECT 1020.580 500.640 1021.700 501.760 ;
 END
END DIB37
PIN DOB37
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1007.560 500.640 1008.680 501.760 ;
  LAYER metal4 ;
  RECT 1007.560 500.640 1008.680 501.760 ;
  LAYER metal3 ;
  RECT 1007.560 500.640 1008.680 501.760 ;
  LAYER metal2 ;
  RECT 1007.560 500.640 1008.680 501.760 ;
  LAYER metal1 ;
  RECT 1007.560 500.640 1008.680 501.760 ;
 END
END DOB37
PIN DIB36
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 993.920 500.640 995.040 501.760 ;
  LAYER metal4 ;
  RECT 993.920 500.640 995.040 501.760 ;
  LAYER metal3 ;
  RECT 993.920 500.640 995.040 501.760 ;
  LAYER metal2 ;
  RECT 993.920 500.640 995.040 501.760 ;
  LAYER metal1 ;
  RECT 993.920 500.640 995.040 501.760 ;
 END
END DIB36
PIN DOB36
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 980.280 500.640 981.400 501.760 ;
  LAYER metal4 ;
  RECT 980.280 500.640 981.400 501.760 ;
  LAYER metal3 ;
  RECT 980.280 500.640 981.400 501.760 ;
  LAYER metal2 ;
  RECT 980.280 500.640 981.400 501.760 ;
  LAYER metal1 ;
  RECT 980.280 500.640 981.400 501.760 ;
 END
END DOB36
PIN DIB35
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 967.260 500.640 968.380 501.760 ;
  LAYER metal4 ;
  RECT 967.260 500.640 968.380 501.760 ;
  LAYER metal3 ;
  RECT 967.260 500.640 968.380 501.760 ;
  LAYER metal2 ;
  RECT 967.260 500.640 968.380 501.760 ;
  LAYER metal1 ;
  RECT 967.260 500.640 968.380 501.760 ;
 END
END DIB35
PIN DOB35
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 953.620 500.640 954.740 501.760 ;
  LAYER metal4 ;
  RECT 953.620 500.640 954.740 501.760 ;
  LAYER metal3 ;
  RECT 953.620 500.640 954.740 501.760 ;
  LAYER metal2 ;
  RECT 953.620 500.640 954.740 501.760 ;
  LAYER metal1 ;
  RECT 953.620 500.640 954.740 501.760 ;
 END
END DOB35
PIN DIB34
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 939.980 500.640 941.100 501.760 ;
  LAYER metal4 ;
  RECT 939.980 500.640 941.100 501.760 ;
  LAYER metal3 ;
  RECT 939.980 500.640 941.100 501.760 ;
  LAYER metal2 ;
  RECT 939.980 500.640 941.100 501.760 ;
  LAYER metal1 ;
  RECT 939.980 500.640 941.100 501.760 ;
 END
END DIB34
PIN DOB34
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 926.960 500.640 928.080 501.760 ;
  LAYER metal4 ;
  RECT 926.960 500.640 928.080 501.760 ;
  LAYER metal3 ;
  RECT 926.960 500.640 928.080 501.760 ;
  LAYER metal2 ;
  RECT 926.960 500.640 928.080 501.760 ;
  LAYER metal1 ;
  RECT 926.960 500.640 928.080 501.760 ;
 END
END DOB34
PIN DIB33
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 913.320 500.640 914.440 501.760 ;
  LAYER metal4 ;
  RECT 913.320 500.640 914.440 501.760 ;
  LAYER metal3 ;
  RECT 913.320 500.640 914.440 501.760 ;
  LAYER metal2 ;
  RECT 913.320 500.640 914.440 501.760 ;
  LAYER metal1 ;
  RECT 913.320 500.640 914.440 501.760 ;
 END
END DIB33
PIN DOB33
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 899.680 500.640 900.800 501.760 ;
  LAYER metal4 ;
  RECT 899.680 500.640 900.800 501.760 ;
  LAYER metal3 ;
  RECT 899.680 500.640 900.800 501.760 ;
  LAYER metal2 ;
  RECT 899.680 500.640 900.800 501.760 ;
  LAYER metal1 ;
  RECT 899.680 500.640 900.800 501.760 ;
 END
END DOB33
PIN DIB32
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 886.040 500.640 887.160 501.760 ;
  LAYER metal4 ;
  RECT 886.040 500.640 887.160 501.760 ;
  LAYER metal3 ;
  RECT 886.040 500.640 887.160 501.760 ;
  LAYER metal2 ;
  RECT 886.040 500.640 887.160 501.760 ;
  LAYER metal1 ;
  RECT 886.040 500.640 887.160 501.760 ;
 END
END DIB32
PIN DOB32
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 873.020 500.640 874.140 501.760 ;
  LAYER metal4 ;
  RECT 873.020 500.640 874.140 501.760 ;
  LAYER metal3 ;
  RECT 873.020 500.640 874.140 501.760 ;
  LAYER metal2 ;
  RECT 873.020 500.640 874.140 501.760 ;
  LAYER metal1 ;
  RECT 873.020 500.640 874.140 501.760 ;
 END
END DOB32
PIN DIB31
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 859.380 500.640 860.500 501.760 ;
  LAYER metal4 ;
  RECT 859.380 500.640 860.500 501.760 ;
  LAYER metal3 ;
  RECT 859.380 500.640 860.500 501.760 ;
  LAYER metal2 ;
  RECT 859.380 500.640 860.500 501.760 ;
  LAYER metal1 ;
  RECT 859.380 500.640 860.500 501.760 ;
 END
END DIB31
PIN DOB31
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 845.740 500.640 846.860 501.760 ;
  LAYER metal4 ;
  RECT 845.740 500.640 846.860 501.760 ;
  LAYER metal3 ;
  RECT 845.740 500.640 846.860 501.760 ;
  LAYER metal2 ;
  RECT 845.740 500.640 846.860 501.760 ;
  LAYER metal1 ;
  RECT 845.740 500.640 846.860 501.760 ;
 END
END DOB31
PIN DIB30
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 832.720 500.640 833.840 501.760 ;
  LAYER metal4 ;
  RECT 832.720 500.640 833.840 501.760 ;
  LAYER metal3 ;
  RECT 832.720 500.640 833.840 501.760 ;
  LAYER metal2 ;
  RECT 832.720 500.640 833.840 501.760 ;
  LAYER metal1 ;
  RECT 832.720 500.640 833.840 501.760 ;
 END
END DIB30
PIN DOB30
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 819.080 500.640 820.200 501.760 ;
  LAYER metal4 ;
  RECT 819.080 500.640 820.200 501.760 ;
  LAYER metal3 ;
  RECT 819.080 500.640 820.200 501.760 ;
  LAYER metal2 ;
  RECT 819.080 500.640 820.200 501.760 ;
  LAYER metal1 ;
  RECT 819.080 500.640 820.200 501.760 ;
 END
END DOB30
PIN DIB29
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 805.440 500.640 806.560 501.760 ;
  LAYER metal4 ;
  RECT 805.440 500.640 806.560 501.760 ;
  LAYER metal3 ;
  RECT 805.440 500.640 806.560 501.760 ;
  LAYER metal2 ;
  RECT 805.440 500.640 806.560 501.760 ;
  LAYER metal1 ;
  RECT 805.440 500.640 806.560 501.760 ;
 END
END DIB29
PIN DOB29
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 792.420 500.640 793.540 501.760 ;
  LAYER metal4 ;
  RECT 792.420 500.640 793.540 501.760 ;
  LAYER metal3 ;
  RECT 792.420 500.640 793.540 501.760 ;
  LAYER metal2 ;
  RECT 792.420 500.640 793.540 501.760 ;
  LAYER metal1 ;
  RECT 792.420 500.640 793.540 501.760 ;
 END
END DOB29
PIN DIB28
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 778.780 500.640 779.900 501.760 ;
  LAYER metal4 ;
  RECT 778.780 500.640 779.900 501.760 ;
  LAYER metal3 ;
  RECT 778.780 500.640 779.900 501.760 ;
  LAYER metal2 ;
  RECT 778.780 500.640 779.900 501.760 ;
  LAYER metal1 ;
  RECT 778.780 500.640 779.900 501.760 ;
 END
END DIB28
PIN DOB28
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 765.140 500.640 766.260 501.760 ;
  LAYER metal4 ;
  RECT 765.140 500.640 766.260 501.760 ;
  LAYER metal3 ;
  RECT 765.140 500.640 766.260 501.760 ;
  LAYER metal2 ;
  RECT 765.140 500.640 766.260 501.760 ;
  LAYER metal1 ;
  RECT 765.140 500.640 766.260 501.760 ;
 END
END DOB28
PIN DIB27
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 752.120 500.640 753.240 501.760 ;
  LAYER metal4 ;
  RECT 752.120 500.640 753.240 501.760 ;
  LAYER metal3 ;
  RECT 752.120 500.640 753.240 501.760 ;
  LAYER metal2 ;
  RECT 752.120 500.640 753.240 501.760 ;
  LAYER metal1 ;
  RECT 752.120 500.640 753.240 501.760 ;
 END
END DIB27
PIN DOB27
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 738.480 500.640 739.600 501.760 ;
  LAYER metal4 ;
  RECT 738.480 500.640 739.600 501.760 ;
  LAYER metal3 ;
  RECT 738.480 500.640 739.600 501.760 ;
  LAYER metal2 ;
  RECT 738.480 500.640 739.600 501.760 ;
  LAYER metal1 ;
  RECT 738.480 500.640 739.600 501.760 ;
 END
END DOB27
PIN DIB26
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 724.840 500.640 725.960 501.760 ;
  LAYER metal4 ;
  RECT 724.840 500.640 725.960 501.760 ;
  LAYER metal3 ;
  RECT 724.840 500.640 725.960 501.760 ;
  LAYER metal2 ;
  RECT 724.840 500.640 725.960 501.760 ;
  LAYER metal1 ;
  RECT 724.840 500.640 725.960 501.760 ;
 END
END DIB26
PIN DOB26
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 711.820 500.640 712.940 501.760 ;
  LAYER metal4 ;
  RECT 711.820 500.640 712.940 501.760 ;
  LAYER metal3 ;
  RECT 711.820 500.640 712.940 501.760 ;
  LAYER metal2 ;
  RECT 711.820 500.640 712.940 501.760 ;
  LAYER metal1 ;
  RECT 711.820 500.640 712.940 501.760 ;
 END
END DOB26
PIN DIB25
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 698.180 500.640 699.300 501.760 ;
  LAYER metal4 ;
  RECT 698.180 500.640 699.300 501.760 ;
  LAYER metal3 ;
  RECT 698.180 500.640 699.300 501.760 ;
  LAYER metal2 ;
  RECT 698.180 500.640 699.300 501.760 ;
  LAYER metal1 ;
  RECT 698.180 500.640 699.300 501.760 ;
 END
END DIB25
PIN DOB25
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 684.540 500.640 685.660 501.760 ;
  LAYER metal4 ;
  RECT 684.540 500.640 685.660 501.760 ;
  LAYER metal3 ;
  RECT 684.540 500.640 685.660 501.760 ;
  LAYER metal2 ;
  RECT 684.540 500.640 685.660 501.760 ;
  LAYER metal1 ;
  RECT 684.540 500.640 685.660 501.760 ;
 END
END DOB25
PIN DIB24
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 671.520 500.640 672.640 501.760 ;
  LAYER metal4 ;
  RECT 671.520 500.640 672.640 501.760 ;
  LAYER metal3 ;
  RECT 671.520 500.640 672.640 501.760 ;
  LAYER metal2 ;
  RECT 671.520 500.640 672.640 501.760 ;
  LAYER metal1 ;
  RECT 671.520 500.640 672.640 501.760 ;
 END
END DIB24
PIN DOB24
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 657.880 500.640 659.000 501.760 ;
  LAYER metal4 ;
  RECT 657.880 500.640 659.000 501.760 ;
  LAYER metal3 ;
  RECT 657.880 500.640 659.000 501.760 ;
  LAYER metal2 ;
  RECT 657.880 500.640 659.000 501.760 ;
  LAYER metal1 ;
  RECT 657.880 500.640 659.000 501.760 ;
 END
END DOB24
PIN DIB23
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 644.240 500.640 645.360 501.760 ;
  LAYER metal4 ;
  RECT 644.240 500.640 645.360 501.760 ;
  LAYER metal3 ;
  RECT 644.240 500.640 645.360 501.760 ;
  LAYER metal2 ;
  RECT 644.240 500.640 645.360 501.760 ;
  LAYER metal1 ;
  RECT 644.240 500.640 645.360 501.760 ;
 END
END DIB23
PIN DOB23
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 631.220 500.640 632.340 501.760 ;
  LAYER metal4 ;
  RECT 631.220 500.640 632.340 501.760 ;
  LAYER metal3 ;
  RECT 631.220 500.640 632.340 501.760 ;
  LAYER metal2 ;
  RECT 631.220 500.640 632.340 501.760 ;
  LAYER metal1 ;
  RECT 631.220 500.640 632.340 501.760 ;
 END
END DOB23
PIN DIB22
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 617.580 500.640 618.700 501.760 ;
  LAYER metal4 ;
  RECT 617.580 500.640 618.700 501.760 ;
  LAYER metal3 ;
  RECT 617.580 500.640 618.700 501.760 ;
  LAYER metal2 ;
  RECT 617.580 500.640 618.700 501.760 ;
  LAYER metal1 ;
  RECT 617.580 500.640 618.700 501.760 ;
 END
END DIB22
PIN DOB22
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 603.940 500.640 605.060 501.760 ;
  LAYER metal4 ;
  RECT 603.940 500.640 605.060 501.760 ;
  LAYER metal3 ;
  RECT 603.940 500.640 605.060 501.760 ;
  LAYER metal2 ;
  RECT 603.940 500.640 605.060 501.760 ;
  LAYER metal1 ;
  RECT 603.940 500.640 605.060 501.760 ;
 END
END DOB22
PIN DIB21
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 590.920 500.640 592.040 501.760 ;
  LAYER metal4 ;
  RECT 590.920 500.640 592.040 501.760 ;
  LAYER metal3 ;
  RECT 590.920 500.640 592.040 501.760 ;
  LAYER metal2 ;
  RECT 590.920 500.640 592.040 501.760 ;
  LAYER metal1 ;
  RECT 590.920 500.640 592.040 501.760 ;
 END
END DIB21
PIN DOB21
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 577.280 500.640 578.400 501.760 ;
  LAYER metal4 ;
  RECT 577.280 500.640 578.400 501.760 ;
  LAYER metal3 ;
  RECT 577.280 500.640 578.400 501.760 ;
  LAYER metal2 ;
  RECT 577.280 500.640 578.400 501.760 ;
  LAYER metal1 ;
  RECT 577.280 500.640 578.400 501.760 ;
 END
END DOB21
PIN DIB20
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 563.640 500.640 564.760 501.760 ;
  LAYER metal4 ;
  RECT 563.640 500.640 564.760 501.760 ;
  LAYER metal3 ;
  RECT 563.640 500.640 564.760 501.760 ;
  LAYER metal2 ;
  RECT 563.640 500.640 564.760 501.760 ;
  LAYER metal1 ;
  RECT 563.640 500.640 564.760 501.760 ;
 END
END DIB20
PIN DOB20
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 550.620 500.640 551.740 501.760 ;
  LAYER metal4 ;
  RECT 550.620 500.640 551.740 501.760 ;
  LAYER metal3 ;
  RECT 550.620 500.640 551.740 501.760 ;
  LAYER metal2 ;
  RECT 550.620 500.640 551.740 501.760 ;
  LAYER metal1 ;
  RECT 550.620 500.640 551.740 501.760 ;
 END
END DOB20
PIN DIB19
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 536.980 500.640 538.100 501.760 ;
  LAYER metal4 ;
  RECT 536.980 500.640 538.100 501.760 ;
  LAYER metal3 ;
  RECT 536.980 500.640 538.100 501.760 ;
  LAYER metal2 ;
  RECT 536.980 500.640 538.100 501.760 ;
  LAYER metal1 ;
  RECT 536.980 500.640 538.100 501.760 ;
 END
END DIB19
PIN DOB19
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 523.340 500.640 524.460 501.760 ;
  LAYER metal4 ;
  RECT 523.340 500.640 524.460 501.760 ;
  LAYER metal3 ;
  RECT 523.340 500.640 524.460 501.760 ;
  LAYER metal2 ;
  RECT 523.340 500.640 524.460 501.760 ;
  LAYER metal1 ;
  RECT 523.340 500.640 524.460 501.760 ;
 END
END DOB19
PIN DIB18
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 510.320 500.640 511.440 501.760 ;
  LAYER metal4 ;
  RECT 510.320 500.640 511.440 501.760 ;
  LAYER metal3 ;
  RECT 510.320 500.640 511.440 501.760 ;
  LAYER metal2 ;
  RECT 510.320 500.640 511.440 501.760 ;
  LAYER metal1 ;
  RECT 510.320 500.640 511.440 501.760 ;
 END
END DIB18
PIN DOB18
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 496.680 500.640 497.800 501.760 ;
  LAYER metal4 ;
  RECT 496.680 500.640 497.800 501.760 ;
  LAYER metal3 ;
  RECT 496.680 500.640 497.800 501.760 ;
  LAYER metal2 ;
  RECT 496.680 500.640 497.800 501.760 ;
  LAYER metal1 ;
  RECT 496.680 500.640 497.800 501.760 ;
 END
END DOB18
PIN DIB17
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 483.040 500.640 484.160 501.760 ;
  LAYER metal4 ;
  RECT 483.040 500.640 484.160 501.760 ;
  LAYER metal3 ;
  RECT 483.040 500.640 484.160 501.760 ;
  LAYER metal2 ;
  RECT 483.040 500.640 484.160 501.760 ;
  LAYER metal1 ;
  RECT 483.040 500.640 484.160 501.760 ;
 END
END DIB17
PIN DOB17
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 469.400 500.640 470.520 501.760 ;
  LAYER metal4 ;
  RECT 469.400 500.640 470.520 501.760 ;
  LAYER metal3 ;
  RECT 469.400 500.640 470.520 501.760 ;
  LAYER metal2 ;
  RECT 469.400 500.640 470.520 501.760 ;
  LAYER metal1 ;
  RECT 469.400 500.640 470.520 501.760 ;
 END
END DOB17
PIN DIB16
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 456.380 500.640 457.500 501.760 ;
  LAYER metal4 ;
  RECT 456.380 500.640 457.500 501.760 ;
  LAYER metal3 ;
  RECT 456.380 500.640 457.500 501.760 ;
  LAYER metal2 ;
  RECT 456.380 500.640 457.500 501.760 ;
  LAYER metal1 ;
  RECT 456.380 500.640 457.500 501.760 ;
 END
END DIB16
PIN DOB16
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 442.740 500.640 443.860 501.760 ;
  LAYER metal4 ;
  RECT 442.740 500.640 443.860 501.760 ;
  LAYER metal3 ;
  RECT 442.740 500.640 443.860 501.760 ;
  LAYER metal2 ;
  RECT 442.740 500.640 443.860 501.760 ;
  LAYER metal1 ;
  RECT 442.740 500.640 443.860 501.760 ;
 END
END DOB16
PIN DIB15
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 429.100 500.640 430.220 501.760 ;
  LAYER metal4 ;
  RECT 429.100 500.640 430.220 501.760 ;
  LAYER metal3 ;
  RECT 429.100 500.640 430.220 501.760 ;
  LAYER metal2 ;
  RECT 429.100 500.640 430.220 501.760 ;
  LAYER metal1 ;
  RECT 429.100 500.640 430.220 501.760 ;
 END
END DIB15
PIN DOB15
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 416.080 500.640 417.200 501.760 ;
  LAYER metal4 ;
  RECT 416.080 500.640 417.200 501.760 ;
  LAYER metal3 ;
  RECT 416.080 500.640 417.200 501.760 ;
  LAYER metal2 ;
  RECT 416.080 500.640 417.200 501.760 ;
  LAYER metal1 ;
  RECT 416.080 500.640 417.200 501.760 ;
 END
END DOB15
PIN DIB14
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 402.440 500.640 403.560 501.760 ;
  LAYER metal4 ;
  RECT 402.440 500.640 403.560 501.760 ;
  LAYER metal3 ;
  RECT 402.440 500.640 403.560 501.760 ;
  LAYER metal2 ;
  RECT 402.440 500.640 403.560 501.760 ;
  LAYER metal1 ;
  RECT 402.440 500.640 403.560 501.760 ;
 END
END DIB14
PIN DOB14
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 388.800 500.640 389.920 501.760 ;
  LAYER metal4 ;
  RECT 388.800 500.640 389.920 501.760 ;
  LAYER metal3 ;
  RECT 388.800 500.640 389.920 501.760 ;
  LAYER metal2 ;
  RECT 388.800 500.640 389.920 501.760 ;
  LAYER metal1 ;
  RECT 388.800 500.640 389.920 501.760 ;
 END
END DOB14
PIN DIB13
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 375.780 500.640 376.900 501.760 ;
  LAYER metal4 ;
  RECT 375.780 500.640 376.900 501.760 ;
  LAYER metal3 ;
  RECT 375.780 500.640 376.900 501.760 ;
  LAYER metal2 ;
  RECT 375.780 500.640 376.900 501.760 ;
  LAYER metal1 ;
  RECT 375.780 500.640 376.900 501.760 ;
 END
END DIB13
PIN DOB13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 362.140 500.640 363.260 501.760 ;
  LAYER metal4 ;
  RECT 362.140 500.640 363.260 501.760 ;
  LAYER metal3 ;
  RECT 362.140 500.640 363.260 501.760 ;
  LAYER metal2 ;
  RECT 362.140 500.640 363.260 501.760 ;
  LAYER metal1 ;
  RECT 362.140 500.640 363.260 501.760 ;
 END
END DOB13
PIN DIB12
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 348.500 500.640 349.620 501.760 ;
  LAYER metal4 ;
  RECT 348.500 500.640 349.620 501.760 ;
  LAYER metal3 ;
  RECT 348.500 500.640 349.620 501.760 ;
  LAYER metal2 ;
  RECT 348.500 500.640 349.620 501.760 ;
  LAYER metal1 ;
  RECT 348.500 500.640 349.620 501.760 ;
 END
END DIB12
PIN DOB12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 335.480 500.640 336.600 501.760 ;
  LAYER metal4 ;
  RECT 335.480 500.640 336.600 501.760 ;
  LAYER metal3 ;
  RECT 335.480 500.640 336.600 501.760 ;
  LAYER metal2 ;
  RECT 335.480 500.640 336.600 501.760 ;
  LAYER metal1 ;
  RECT 335.480 500.640 336.600 501.760 ;
 END
END DOB12
PIN DIB11
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 321.840 500.640 322.960 501.760 ;
  LAYER metal4 ;
  RECT 321.840 500.640 322.960 501.760 ;
  LAYER metal3 ;
  RECT 321.840 500.640 322.960 501.760 ;
  LAYER metal2 ;
  RECT 321.840 500.640 322.960 501.760 ;
  LAYER metal1 ;
  RECT 321.840 500.640 322.960 501.760 ;
 END
END DIB11
PIN DOB11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 308.200 500.640 309.320 501.760 ;
  LAYER metal4 ;
  RECT 308.200 500.640 309.320 501.760 ;
  LAYER metal3 ;
  RECT 308.200 500.640 309.320 501.760 ;
  LAYER metal2 ;
  RECT 308.200 500.640 309.320 501.760 ;
  LAYER metal1 ;
  RECT 308.200 500.640 309.320 501.760 ;
 END
END DOB11
PIN DIB10
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 295.180 500.640 296.300 501.760 ;
  LAYER metal4 ;
  RECT 295.180 500.640 296.300 501.760 ;
  LAYER metal3 ;
  RECT 295.180 500.640 296.300 501.760 ;
  LAYER metal2 ;
  RECT 295.180 500.640 296.300 501.760 ;
  LAYER metal1 ;
  RECT 295.180 500.640 296.300 501.760 ;
 END
END DIB10
PIN DOB10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 281.540 500.640 282.660 501.760 ;
  LAYER metal4 ;
  RECT 281.540 500.640 282.660 501.760 ;
  LAYER metal3 ;
  RECT 281.540 500.640 282.660 501.760 ;
  LAYER metal2 ;
  RECT 281.540 500.640 282.660 501.760 ;
  LAYER metal1 ;
  RECT 281.540 500.640 282.660 501.760 ;
 END
END DOB10
PIN DIB9
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 267.900 500.640 269.020 501.760 ;
  LAYER metal4 ;
  RECT 267.900 500.640 269.020 501.760 ;
  LAYER metal3 ;
  RECT 267.900 500.640 269.020 501.760 ;
  LAYER metal2 ;
  RECT 267.900 500.640 269.020 501.760 ;
  LAYER metal1 ;
  RECT 267.900 500.640 269.020 501.760 ;
 END
END DIB9
PIN DOB9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 254.880 500.640 256.000 501.760 ;
  LAYER metal4 ;
  RECT 254.880 500.640 256.000 501.760 ;
  LAYER metal3 ;
  RECT 254.880 500.640 256.000 501.760 ;
  LAYER metal2 ;
  RECT 254.880 500.640 256.000 501.760 ;
  LAYER metal1 ;
  RECT 254.880 500.640 256.000 501.760 ;
 END
END DOB9
PIN DIB8
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 241.240 500.640 242.360 501.760 ;
  LAYER metal4 ;
  RECT 241.240 500.640 242.360 501.760 ;
  LAYER metal3 ;
  RECT 241.240 500.640 242.360 501.760 ;
  LAYER metal2 ;
  RECT 241.240 500.640 242.360 501.760 ;
  LAYER metal1 ;
  RECT 241.240 500.640 242.360 501.760 ;
 END
END DIB8
PIN DOB8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 227.600 500.640 228.720 501.760 ;
  LAYER metal4 ;
  RECT 227.600 500.640 228.720 501.760 ;
  LAYER metal3 ;
  RECT 227.600 500.640 228.720 501.760 ;
  LAYER metal2 ;
  RECT 227.600 500.640 228.720 501.760 ;
  LAYER metal1 ;
  RECT 227.600 500.640 228.720 501.760 ;
 END
END DOB8
PIN DIB7
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 214.580 500.640 215.700 501.760 ;
  LAYER metal4 ;
  RECT 214.580 500.640 215.700 501.760 ;
  LAYER metal3 ;
  RECT 214.580 500.640 215.700 501.760 ;
  LAYER metal2 ;
  RECT 214.580 500.640 215.700 501.760 ;
  LAYER metal1 ;
  RECT 214.580 500.640 215.700 501.760 ;
 END
END DIB7
PIN DOB7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 200.940 500.640 202.060 501.760 ;
  LAYER metal4 ;
  RECT 200.940 500.640 202.060 501.760 ;
  LAYER metal3 ;
  RECT 200.940 500.640 202.060 501.760 ;
  LAYER metal2 ;
  RECT 200.940 500.640 202.060 501.760 ;
  LAYER metal1 ;
  RECT 200.940 500.640 202.060 501.760 ;
 END
END DOB7
PIN DIB6
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 187.300 500.640 188.420 501.760 ;
  LAYER metal4 ;
  RECT 187.300 500.640 188.420 501.760 ;
  LAYER metal3 ;
  RECT 187.300 500.640 188.420 501.760 ;
  LAYER metal2 ;
  RECT 187.300 500.640 188.420 501.760 ;
  LAYER metal1 ;
  RECT 187.300 500.640 188.420 501.760 ;
 END
END DIB6
PIN DOB6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 174.280 500.640 175.400 501.760 ;
  LAYER metal4 ;
  RECT 174.280 500.640 175.400 501.760 ;
  LAYER metal3 ;
  RECT 174.280 500.640 175.400 501.760 ;
  LAYER metal2 ;
  RECT 174.280 500.640 175.400 501.760 ;
  LAYER metal1 ;
  RECT 174.280 500.640 175.400 501.760 ;
 END
END DOB6
PIN DIB5
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 160.640 500.640 161.760 501.760 ;
  LAYER metal4 ;
  RECT 160.640 500.640 161.760 501.760 ;
  LAYER metal3 ;
  RECT 160.640 500.640 161.760 501.760 ;
  LAYER metal2 ;
  RECT 160.640 500.640 161.760 501.760 ;
  LAYER metal1 ;
  RECT 160.640 500.640 161.760 501.760 ;
 END
END DIB5
PIN DOB5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 147.000 500.640 148.120 501.760 ;
  LAYER metal4 ;
  RECT 147.000 500.640 148.120 501.760 ;
  LAYER metal3 ;
  RECT 147.000 500.640 148.120 501.760 ;
  LAYER metal2 ;
  RECT 147.000 500.640 148.120 501.760 ;
  LAYER metal1 ;
  RECT 147.000 500.640 148.120 501.760 ;
 END
END DOB5
PIN DIB4
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 133.980 500.640 135.100 501.760 ;
  LAYER metal4 ;
  RECT 133.980 500.640 135.100 501.760 ;
  LAYER metal3 ;
  RECT 133.980 500.640 135.100 501.760 ;
  LAYER metal2 ;
  RECT 133.980 500.640 135.100 501.760 ;
  LAYER metal1 ;
  RECT 133.980 500.640 135.100 501.760 ;
 END
END DIB4
PIN DOB4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 120.340 500.640 121.460 501.760 ;
  LAYER metal4 ;
  RECT 120.340 500.640 121.460 501.760 ;
  LAYER metal3 ;
  RECT 120.340 500.640 121.460 501.760 ;
  LAYER metal2 ;
  RECT 120.340 500.640 121.460 501.760 ;
  LAYER metal1 ;
  RECT 120.340 500.640 121.460 501.760 ;
 END
END DOB4
PIN DIB3
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 106.700 500.640 107.820 501.760 ;
  LAYER metal4 ;
  RECT 106.700 500.640 107.820 501.760 ;
  LAYER metal3 ;
  RECT 106.700 500.640 107.820 501.760 ;
  LAYER metal2 ;
  RECT 106.700 500.640 107.820 501.760 ;
  LAYER metal1 ;
  RECT 106.700 500.640 107.820 501.760 ;
 END
END DIB3
PIN DOB3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 93.680 500.640 94.800 501.760 ;
  LAYER metal4 ;
  RECT 93.680 500.640 94.800 501.760 ;
  LAYER metal3 ;
  RECT 93.680 500.640 94.800 501.760 ;
  LAYER metal2 ;
  RECT 93.680 500.640 94.800 501.760 ;
  LAYER metal1 ;
  RECT 93.680 500.640 94.800 501.760 ;
 END
END DOB3
PIN DIB2
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 80.040 500.640 81.160 501.760 ;
  LAYER metal4 ;
  RECT 80.040 500.640 81.160 501.760 ;
  LAYER metal3 ;
  RECT 80.040 500.640 81.160 501.760 ;
  LAYER metal2 ;
  RECT 80.040 500.640 81.160 501.760 ;
  LAYER metal1 ;
  RECT 80.040 500.640 81.160 501.760 ;
 END
END DIB2
PIN DOB2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 66.400 500.640 67.520 501.760 ;
  LAYER metal4 ;
  RECT 66.400 500.640 67.520 501.760 ;
  LAYER metal3 ;
  RECT 66.400 500.640 67.520 501.760 ;
  LAYER metal2 ;
  RECT 66.400 500.640 67.520 501.760 ;
  LAYER metal1 ;
  RECT 66.400 500.640 67.520 501.760 ;
 END
END DOB2
PIN DIB1
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 52.760 500.640 53.880 501.760 ;
  LAYER metal4 ;
  RECT 52.760 500.640 53.880 501.760 ;
  LAYER metal3 ;
  RECT 52.760 500.640 53.880 501.760 ;
  LAYER metal2 ;
  RECT 52.760 500.640 53.880 501.760 ;
  LAYER metal1 ;
  RECT 52.760 500.640 53.880 501.760 ;
 END
END DIB1
PIN DOB1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 39.740 500.640 40.860 501.760 ;
  LAYER metal4 ;
  RECT 39.740 500.640 40.860 501.760 ;
  LAYER metal3 ;
  RECT 39.740 500.640 40.860 501.760 ;
  LAYER metal2 ;
  RECT 39.740 500.640 40.860 501.760 ;
  LAYER metal1 ;
  RECT 39.740 500.640 40.860 501.760 ;
 END
END DOB1
PIN DIB0
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 26.100 500.640 27.220 501.760 ;
  LAYER metal4 ;
  RECT 26.100 500.640 27.220 501.760 ;
  LAYER metal3 ;
  RECT 26.100 500.640 27.220 501.760 ;
  LAYER metal2 ;
  RECT 26.100 500.640 27.220 501.760 ;
  LAYER metal1 ;
  RECT 26.100 500.640 27.220 501.760 ;
 END
END DIB0
PIN DOB0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 12.460 500.640 13.580 501.760 ;
  LAYER metal4 ;
  RECT 12.460 500.640 13.580 501.760 ;
  LAYER metal3 ;
  RECT 12.460 500.640 13.580 501.760 ;
  LAYER metal2 ;
  RECT 12.460 500.640 13.580 501.760 ;
  LAYER metal1 ;
  RECT 12.460 500.640 13.580 501.760 ;
 END
END DOB0
PIN DIA127
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3573.120 0.000 3574.240 1.120 ;
  LAYER metal4 ;
  RECT 3573.120 0.000 3574.240 1.120 ;
  LAYER metal3 ;
  RECT 3573.120 0.000 3574.240 1.120 ;
  LAYER metal2 ;
  RECT 3573.120 0.000 3574.240 1.120 ;
  LAYER metal1 ;
  RECT 3573.120 0.000 3574.240 1.120 ;
 END
END DIA127
PIN DOA127
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3559.480 0.000 3560.600 1.120 ;
  LAYER metal4 ;
  RECT 3559.480 0.000 3560.600 1.120 ;
  LAYER metal3 ;
  RECT 3559.480 0.000 3560.600 1.120 ;
  LAYER metal2 ;
  RECT 3559.480 0.000 3560.600 1.120 ;
  LAYER metal1 ;
  RECT 3559.480 0.000 3560.600 1.120 ;
 END
END DOA127
PIN DIA126
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3546.460 0.000 3547.580 1.120 ;
  LAYER metal4 ;
  RECT 3546.460 0.000 3547.580 1.120 ;
  LAYER metal3 ;
  RECT 3546.460 0.000 3547.580 1.120 ;
  LAYER metal2 ;
  RECT 3546.460 0.000 3547.580 1.120 ;
  LAYER metal1 ;
  RECT 3546.460 0.000 3547.580 1.120 ;
 END
END DIA126
PIN DOA126
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3532.820 0.000 3533.940 1.120 ;
  LAYER metal4 ;
  RECT 3532.820 0.000 3533.940 1.120 ;
  LAYER metal3 ;
  RECT 3532.820 0.000 3533.940 1.120 ;
  LAYER metal2 ;
  RECT 3532.820 0.000 3533.940 1.120 ;
  LAYER metal1 ;
  RECT 3532.820 0.000 3533.940 1.120 ;
 END
END DOA126
PIN DIA125
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3519.180 0.000 3520.300 1.120 ;
  LAYER metal4 ;
  RECT 3519.180 0.000 3520.300 1.120 ;
  LAYER metal3 ;
  RECT 3519.180 0.000 3520.300 1.120 ;
  LAYER metal2 ;
  RECT 3519.180 0.000 3520.300 1.120 ;
  LAYER metal1 ;
  RECT 3519.180 0.000 3520.300 1.120 ;
 END
END DIA125
PIN DOA125
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3506.160 0.000 3507.280 1.120 ;
  LAYER metal4 ;
  RECT 3506.160 0.000 3507.280 1.120 ;
  LAYER metal3 ;
  RECT 3506.160 0.000 3507.280 1.120 ;
  LAYER metal2 ;
  RECT 3506.160 0.000 3507.280 1.120 ;
  LAYER metal1 ;
  RECT 3506.160 0.000 3507.280 1.120 ;
 END
END DOA125
PIN DIA124
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3492.520 0.000 3493.640 1.120 ;
  LAYER metal4 ;
  RECT 3492.520 0.000 3493.640 1.120 ;
  LAYER metal3 ;
  RECT 3492.520 0.000 3493.640 1.120 ;
  LAYER metal2 ;
  RECT 3492.520 0.000 3493.640 1.120 ;
  LAYER metal1 ;
  RECT 3492.520 0.000 3493.640 1.120 ;
 END
END DIA124
PIN DOA124
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3478.880 0.000 3480.000 1.120 ;
  LAYER metal4 ;
  RECT 3478.880 0.000 3480.000 1.120 ;
  LAYER metal3 ;
  RECT 3478.880 0.000 3480.000 1.120 ;
  LAYER metal2 ;
  RECT 3478.880 0.000 3480.000 1.120 ;
  LAYER metal1 ;
  RECT 3478.880 0.000 3480.000 1.120 ;
 END
END DOA124
PIN DIA123
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3465.860 0.000 3466.980 1.120 ;
  LAYER metal4 ;
  RECT 3465.860 0.000 3466.980 1.120 ;
  LAYER metal3 ;
  RECT 3465.860 0.000 3466.980 1.120 ;
  LAYER metal2 ;
  RECT 3465.860 0.000 3466.980 1.120 ;
  LAYER metal1 ;
  RECT 3465.860 0.000 3466.980 1.120 ;
 END
END DIA123
PIN DOA123
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3452.220 0.000 3453.340 1.120 ;
  LAYER metal4 ;
  RECT 3452.220 0.000 3453.340 1.120 ;
  LAYER metal3 ;
  RECT 3452.220 0.000 3453.340 1.120 ;
  LAYER metal2 ;
  RECT 3452.220 0.000 3453.340 1.120 ;
  LAYER metal1 ;
  RECT 3452.220 0.000 3453.340 1.120 ;
 END
END DOA123
PIN DIA122
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3438.580 0.000 3439.700 1.120 ;
  LAYER metal4 ;
  RECT 3438.580 0.000 3439.700 1.120 ;
  LAYER metal3 ;
  RECT 3438.580 0.000 3439.700 1.120 ;
  LAYER metal2 ;
  RECT 3438.580 0.000 3439.700 1.120 ;
  LAYER metal1 ;
  RECT 3438.580 0.000 3439.700 1.120 ;
 END
END DIA122
PIN DOA122
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3425.560 0.000 3426.680 1.120 ;
  LAYER metal4 ;
  RECT 3425.560 0.000 3426.680 1.120 ;
  LAYER metal3 ;
  RECT 3425.560 0.000 3426.680 1.120 ;
  LAYER metal2 ;
  RECT 3425.560 0.000 3426.680 1.120 ;
  LAYER metal1 ;
  RECT 3425.560 0.000 3426.680 1.120 ;
 END
END DOA122
PIN DIA121
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3411.920 0.000 3413.040 1.120 ;
  LAYER metal4 ;
  RECT 3411.920 0.000 3413.040 1.120 ;
  LAYER metal3 ;
  RECT 3411.920 0.000 3413.040 1.120 ;
  LAYER metal2 ;
  RECT 3411.920 0.000 3413.040 1.120 ;
  LAYER metal1 ;
  RECT 3411.920 0.000 3413.040 1.120 ;
 END
END DIA121
PIN DOA121
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3398.280 0.000 3399.400 1.120 ;
  LAYER metal4 ;
  RECT 3398.280 0.000 3399.400 1.120 ;
  LAYER metal3 ;
  RECT 3398.280 0.000 3399.400 1.120 ;
  LAYER metal2 ;
  RECT 3398.280 0.000 3399.400 1.120 ;
  LAYER metal1 ;
  RECT 3398.280 0.000 3399.400 1.120 ;
 END
END DOA121
PIN DIA120
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3385.260 0.000 3386.380 1.120 ;
  LAYER metal4 ;
  RECT 3385.260 0.000 3386.380 1.120 ;
  LAYER metal3 ;
  RECT 3385.260 0.000 3386.380 1.120 ;
  LAYER metal2 ;
  RECT 3385.260 0.000 3386.380 1.120 ;
  LAYER metal1 ;
  RECT 3385.260 0.000 3386.380 1.120 ;
 END
END DIA120
PIN DOA120
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3371.620 0.000 3372.740 1.120 ;
  LAYER metal4 ;
  RECT 3371.620 0.000 3372.740 1.120 ;
  LAYER metal3 ;
  RECT 3371.620 0.000 3372.740 1.120 ;
  LAYER metal2 ;
  RECT 3371.620 0.000 3372.740 1.120 ;
  LAYER metal1 ;
  RECT 3371.620 0.000 3372.740 1.120 ;
 END
END DOA120
PIN DIA119
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3357.980 0.000 3359.100 1.120 ;
  LAYER metal4 ;
  RECT 3357.980 0.000 3359.100 1.120 ;
  LAYER metal3 ;
  RECT 3357.980 0.000 3359.100 1.120 ;
  LAYER metal2 ;
  RECT 3357.980 0.000 3359.100 1.120 ;
  LAYER metal1 ;
  RECT 3357.980 0.000 3359.100 1.120 ;
 END
END DIA119
PIN DOA119
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3344.960 0.000 3346.080 1.120 ;
  LAYER metal4 ;
  RECT 3344.960 0.000 3346.080 1.120 ;
  LAYER metal3 ;
  RECT 3344.960 0.000 3346.080 1.120 ;
  LAYER metal2 ;
  RECT 3344.960 0.000 3346.080 1.120 ;
  LAYER metal1 ;
  RECT 3344.960 0.000 3346.080 1.120 ;
 END
END DOA119
PIN DIA118
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3331.320 0.000 3332.440 1.120 ;
  LAYER metal4 ;
  RECT 3331.320 0.000 3332.440 1.120 ;
  LAYER metal3 ;
  RECT 3331.320 0.000 3332.440 1.120 ;
  LAYER metal2 ;
  RECT 3331.320 0.000 3332.440 1.120 ;
  LAYER metal1 ;
  RECT 3331.320 0.000 3332.440 1.120 ;
 END
END DIA118
PIN DOA118
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3317.680 0.000 3318.800 1.120 ;
  LAYER metal4 ;
  RECT 3317.680 0.000 3318.800 1.120 ;
  LAYER metal3 ;
  RECT 3317.680 0.000 3318.800 1.120 ;
  LAYER metal2 ;
  RECT 3317.680 0.000 3318.800 1.120 ;
  LAYER metal1 ;
  RECT 3317.680 0.000 3318.800 1.120 ;
 END
END DOA118
PIN DIA117
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3304.660 0.000 3305.780 1.120 ;
  LAYER metal4 ;
  RECT 3304.660 0.000 3305.780 1.120 ;
  LAYER metal3 ;
  RECT 3304.660 0.000 3305.780 1.120 ;
  LAYER metal2 ;
  RECT 3304.660 0.000 3305.780 1.120 ;
  LAYER metal1 ;
  RECT 3304.660 0.000 3305.780 1.120 ;
 END
END DIA117
PIN DOA117
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3291.020 0.000 3292.140 1.120 ;
  LAYER metal4 ;
  RECT 3291.020 0.000 3292.140 1.120 ;
  LAYER metal3 ;
  RECT 3291.020 0.000 3292.140 1.120 ;
  LAYER metal2 ;
  RECT 3291.020 0.000 3292.140 1.120 ;
  LAYER metal1 ;
  RECT 3291.020 0.000 3292.140 1.120 ;
 END
END DOA117
PIN DIA116
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3277.380 0.000 3278.500 1.120 ;
  LAYER metal4 ;
  RECT 3277.380 0.000 3278.500 1.120 ;
  LAYER metal3 ;
  RECT 3277.380 0.000 3278.500 1.120 ;
  LAYER metal2 ;
  RECT 3277.380 0.000 3278.500 1.120 ;
  LAYER metal1 ;
  RECT 3277.380 0.000 3278.500 1.120 ;
 END
END DIA116
PIN DOA116
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3264.360 0.000 3265.480 1.120 ;
  LAYER metal4 ;
  RECT 3264.360 0.000 3265.480 1.120 ;
  LAYER metal3 ;
  RECT 3264.360 0.000 3265.480 1.120 ;
  LAYER metal2 ;
  RECT 3264.360 0.000 3265.480 1.120 ;
  LAYER metal1 ;
  RECT 3264.360 0.000 3265.480 1.120 ;
 END
END DOA116
PIN DIA115
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3250.720 0.000 3251.840 1.120 ;
  LAYER metal4 ;
  RECT 3250.720 0.000 3251.840 1.120 ;
  LAYER metal3 ;
  RECT 3250.720 0.000 3251.840 1.120 ;
  LAYER metal2 ;
  RECT 3250.720 0.000 3251.840 1.120 ;
  LAYER metal1 ;
  RECT 3250.720 0.000 3251.840 1.120 ;
 END
END DIA115
PIN DOA115
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3237.080 0.000 3238.200 1.120 ;
  LAYER metal4 ;
  RECT 3237.080 0.000 3238.200 1.120 ;
  LAYER metal3 ;
  RECT 3237.080 0.000 3238.200 1.120 ;
  LAYER metal2 ;
  RECT 3237.080 0.000 3238.200 1.120 ;
  LAYER metal1 ;
  RECT 3237.080 0.000 3238.200 1.120 ;
 END
END DOA115
PIN DIA114
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3224.060 0.000 3225.180 1.120 ;
  LAYER metal4 ;
  RECT 3224.060 0.000 3225.180 1.120 ;
  LAYER metal3 ;
  RECT 3224.060 0.000 3225.180 1.120 ;
  LAYER metal2 ;
  RECT 3224.060 0.000 3225.180 1.120 ;
  LAYER metal1 ;
  RECT 3224.060 0.000 3225.180 1.120 ;
 END
END DIA114
PIN DOA114
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3210.420 0.000 3211.540 1.120 ;
  LAYER metal4 ;
  RECT 3210.420 0.000 3211.540 1.120 ;
  LAYER metal3 ;
  RECT 3210.420 0.000 3211.540 1.120 ;
  LAYER metal2 ;
  RECT 3210.420 0.000 3211.540 1.120 ;
  LAYER metal1 ;
  RECT 3210.420 0.000 3211.540 1.120 ;
 END
END DOA114
PIN DIA113
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3196.780 0.000 3197.900 1.120 ;
  LAYER metal4 ;
  RECT 3196.780 0.000 3197.900 1.120 ;
  LAYER metal3 ;
  RECT 3196.780 0.000 3197.900 1.120 ;
  LAYER metal2 ;
  RECT 3196.780 0.000 3197.900 1.120 ;
  LAYER metal1 ;
  RECT 3196.780 0.000 3197.900 1.120 ;
 END
END DIA113
PIN DOA113
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3183.760 0.000 3184.880 1.120 ;
  LAYER metal4 ;
  RECT 3183.760 0.000 3184.880 1.120 ;
  LAYER metal3 ;
  RECT 3183.760 0.000 3184.880 1.120 ;
  LAYER metal2 ;
  RECT 3183.760 0.000 3184.880 1.120 ;
  LAYER metal1 ;
  RECT 3183.760 0.000 3184.880 1.120 ;
 END
END DOA113
PIN DIA112
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3170.120 0.000 3171.240 1.120 ;
  LAYER metal4 ;
  RECT 3170.120 0.000 3171.240 1.120 ;
  LAYER metal3 ;
  RECT 3170.120 0.000 3171.240 1.120 ;
  LAYER metal2 ;
  RECT 3170.120 0.000 3171.240 1.120 ;
  LAYER metal1 ;
  RECT 3170.120 0.000 3171.240 1.120 ;
 END
END DIA112
PIN DOA112
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3156.480 0.000 3157.600 1.120 ;
  LAYER metal4 ;
  RECT 3156.480 0.000 3157.600 1.120 ;
  LAYER metal3 ;
  RECT 3156.480 0.000 3157.600 1.120 ;
  LAYER metal2 ;
  RECT 3156.480 0.000 3157.600 1.120 ;
  LAYER metal1 ;
  RECT 3156.480 0.000 3157.600 1.120 ;
 END
END DOA112
PIN DIA111
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3142.840 0.000 3143.960 1.120 ;
  LAYER metal4 ;
  RECT 3142.840 0.000 3143.960 1.120 ;
  LAYER metal3 ;
  RECT 3142.840 0.000 3143.960 1.120 ;
  LAYER metal2 ;
  RECT 3142.840 0.000 3143.960 1.120 ;
  LAYER metal1 ;
  RECT 3142.840 0.000 3143.960 1.120 ;
 END
END DIA111
PIN DOA111
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3129.820 0.000 3130.940 1.120 ;
  LAYER metal4 ;
  RECT 3129.820 0.000 3130.940 1.120 ;
  LAYER metal3 ;
  RECT 3129.820 0.000 3130.940 1.120 ;
  LAYER metal2 ;
  RECT 3129.820 0.000 3130.940 1.120 ;
  LAYER metal1 ;
  RECT 3129.820 0.000 3130.940 1.120 ;
 END
END DOA111
PIN DIA110
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3116.180 0.000 3117.300 1.120 ;
  LAYER metal4 ;
  RECT 3116.180 0.000 3117.300 1.120 ;
  LAYER metal3 ;
  RECT 3116.180 0.000 3117.300 1.120 ;
  LAYER metal2 ;
  RECT 3116.180 0.000 3117.300 1.120 ;
  LAYER metal1 ;
  RECT 3116.180 0.000 3117.300 1.120 ;
 END
END DIA110
PIN DOA110
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3102.540 0.000 3103.660 1.120 ;
  LAYER metal4 ;
  RECT 3102.540 0.000 3103.660 1.120 ;
  LAYER metal3 ;
  RECT 3102.540 0.000 3103.660 1.120 ;
  LAYER metal2 ;
  RECT 3102.540 0.000 3103.660 1.120 ;
  LAYER metal1 ;
  RECT 3102.540 0.000 3103.660 1.120 ;
 END
END DOA110
PIN DIA109
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3089.520 0.000 3090.640 1.120 ;
  LAYER metal4 ;
  RECT 3089.520 0.000 3090.640 1.120 ;
  LAYER metal3 ;
  RECT 3089.520 0.000 3090.640 1.120 ;
  LAYER metal2 ;
  RECT 3089.520 0.000 3090.640 1.120 ;
  LAYER metal1 ;
  RECT 3089.520 0.000 3090.640 1.120 ;
 END
END DIA109
PIN DOA109
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3075.880 0.000 3077.000 1.120 ;
  LAYER metal4 ;
  RECT 3075.880 0.000 3077.000 1.120 ;
  LAYER metal3 ;
  RECT 3075.880 0.000 3077.000 1.120 ;
  LAYER metal2 ;
  RECT 3075.880 0.000 3077.000 1.120 ;
  LAYER metal1 ;
  RECT 3075.880 0.000 3077.000 1.120 ;
 END
END DOA109
PIN DIA108
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3062.240 0.000 3063.360 1.120 ;
  LAYER metal4 ;
  RECT 3062.240 0.000 3063.360 1.120 ;
  LAYER metal3 ;
  RECT 3062.240 0.000 3063.360 1.120 ;
  LAYER metal2 ;
  RECT 3062.240 0.000 3063.360 1.120 ;
  LAYER metal1 ;
  RECT 3062.240 0.000 3063.360 1.120 ;
 END
END DIA108
PIN DOA108
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3049.220 0.000 3050.340 1.120 ;
  LAYER metal4 ;
  RECT 3049.220 0.000 3050.340 1.120 ;
  LAYER metal3 ;
  RECT 3049.220 0.000 3050.340 1.120 ;
  LAYER metal2 ;
  RECT 3049.220 0.000 3050.340 1.120 ;
  LAYER metal1 ;
  RECT 3049.220 0.000 3050.340 1.120 ;
 END
END DOA108
PIN DIA107
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3035.580 0.000 3036.700 1.120 ;
  LAYER metal4 ;
  RECT 3035.580 0.000 3036.700 1.120 ;
  LAYER metal3 ;
  RECT 3035.580 0.000 3036.700 1.120 ;
  LAYER metal2 ;
  RECT 3035.580 0.000 3036.700 1.120 ;
  LAYER metal1 ;
  RECT 3035.580 0.000 3036.700 1.120 ;
 END
END DIA107
PIN DOA107
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3021.940 0.000 3023.060 1.120 ;
  LAYER metal4 ;
  RECT 3021.940 0.000 3023.060 1.120 ;
  LAYER metal3 ;
  RECT 3021.940 0.000 3023.060 1.120 ;
  LAYER metal2 ;
  RECT 3021.940 0.000 3023.060 1.120 ;
  LAYER metal1 ;
  RECT 3021.940 0.000 3023.060 1.120 ;
 END
END DOA107
PIN DIA106
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3008.920 0.000 3010.040 1.120 ;
  LAYER metal4 ;
  RECT 3008.920 0.000 3010.040 1.120 ;
  LAYER metal3 ;
  RECT 3008.920 0.000 3010.040 1.120 ;
  LAYER metal2 ;
  RECT 3008.920 0.000 3010.040 1.120 ;
  LAYER metal1 ;
  RECT 3008.920 0.000 3010.040 1.120 ;
 END
END DIA106
PIN DOA106
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2995.280 0.000 2996.400 1.120 ;
  LAYER metal4 ;
  RECT 2995.280 0.000 2996.400 1.120 ;
  LAYER metal3 ;
  RECT 2995.280 0.000 2996.400 1.120 ;
  LAYER metal2 ;
  RECT 2995.280 0.000 2996.400 1.120 ;
  LAYER metal1 ;
  RECT 2995.280 0.000 2996.400 1.120 ;
 END
END DOA106
PIN DIA105
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2981.640 0.000 2982.760 1.120 ;
  LAYER metal4 ;
  RECT 2981.640 0.000 2982.760 1.120 ;
  LAYER metal3 ;
  RECT 2981.640 0.000 2982.760 1.120 ;
  LAYER metal2 ;
  RECT 2981.640 0.000 2982.760 1.120 ;
  LAYER metal1 ;
  RECT 2981.640 0.000 2982.760 1.120 ;
 END
END DIA105
PIN DOA105
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2968.620 0.000 2969.740 1.120 ;
  LAYER metal4 ;
  RECT 2968.620 0.000 2969.740 1.120 ;
  LAYER metal3 ;
  RECT 2968.620 0.000 2969.740 1.120 ;
  LAYER metal2 ;
  RECT 2968.620 0.000 2969.740 1.120 ;
  LAYER metal1 ;
  RECT 2968.620 0.000 2969.740 1.120 ;
 END
END DOA105
PIN DIA104
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2954.980 0.000 2956.100 1.120 ;
  LAYER metal4 ;
  RECT 2954.980 0.000 2956.100 1.120 ;
  LAYER metal3 ;
  RECT 2954.980 0.000 2956.100 1.120 ;
  LAYER metal2 ;
  RECT 2954.980 0.000 2956.100 1.120 ;
  LAYER metal1 ;
  RECT 2954.980 0.000 2956.100 1.120 ;
 END
END DIA104
PIN DOA104
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2941.340 0.000 2942.460 1.120 ;
  LAYER metal4 ;
  RECT 2941.340 0.000 2942.460 1.120 ;
  LAYER metal3 ;
  RECT 2941.340 0.000 2942.460 1.120 ;
  LAYER metal2 ;
  RECT 2941.340 0.000 2942.460 1.120 ;
  LAYER metal1 ;
  RECT 2941.340 0.000 2942.460 1.120 ;
 END
END DOA104
PIN DIA103
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2928.320 0.000 2929.440 1.120 ;
  LAYER metal4 ;
  RECT 2928.320 0.000 2929.440 1.120 ;
  LAYER metal3 ;
  RECT 2928.320 0.000 2929.440 1.120 ;
  LAYER metal2 ;
  RECT 2928.320 0.000 2929.440 1.120 ;
  LAYER metal1 ;
  RECT 2928.320 0.000 2929.440 1.120 ;
 END
END DIA103
PIN DOA103
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2914.680 0.000 2915.800 1.120 ;
  LAYER metal4 ;
  RECT 2914.680 0.000 2915.800 1.120 ;
  LAYER metal3 ;
  RECT 2914.680 0.000 2915.800 1.120 ;
  LAYER metal2 ;
  RECT 2914.680 0.000 2915.800 1.120 ;
  LAYER metal1 ;
  RECT 2914.680 0.000 2915.800 1.120 ;
 END
END DOA103
PIN DIA102
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2901.040 0.000 2902.160 1.120 ;
  LAYER metal4 ;
  RECT 2901.040 0.000 2902.160 1.120 ;
  LAYER metal3 ;
  RECT 2901.040 0.000 2902.160 1.120 ;
  LAYER metal2 ;
  RECT 2901.040 0.000 2902.160 1.120 ;
  LAYER metal1 ;
  RECT 2901.040 0.000 2902.160 1.120 ;
 END
END DIA102
PIN DOA102
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2888.020 0.000 2889.140 1.120 ;
  LAYER metal4 ;
  RECT 2888.020 0.000 2889.140 1.120 ;
  LAYER metal3 ;
  RECT 2888.020 0.000 2889.140 1.120 ;
  LAYER metal2 ;
  RECT 2888.020 0.000 2889.140 1.120 ;
  LAYER metal1 ;
  RECT 2888.020 0.000 2889.140 1.120 ;
 END
END DOA102
PIN DIA101
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2874.380 0.000 2875.500 1.120 ;
  LAYER metal4 ;
  RECT 2874.380 0.000 2875.500 1.120 ;
  LAYER metal3 ;
  RECT 2874.380 0.000 2875.500 1.120 ;
  LAYER metal2 ;
  RECT 2874.380 0.000 2875.500 1.120 ;
  LAYER metal1 ;
  RECT 2874.380 0.000 2875.500 1.120 ;
 END
END DIA101
PIN DOA101
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2860.740 0.000 2861.860 1.120 ;
  LAYER metal4 ;
  RECT 2860.740 0.000 2861.860 1.120 ;
  LAYER metal3 ;
  RECT 2860.740 0.000 2861.860 1.120 ;
  LAYER metal2 ;
  RECT 2860.740 0.000 2861.860 1.120 ;
  LAYER metal1 ;
  RECT 2860.740 0.000 2861.860 1.120 ;
 END
END DOA101
PIN DIA100
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2847.720 0.000 2848.840 1.120 ;
  LAYER metal4 ;
  RECT 2847.720 0.000 2848.840 1.120 ;
  LAYER metal3 ;
  RECT 2847.720 0.000 2848.840 1.120 ;
  LAYER metal2 ;
  RECT 2847.720 0.000 2848.840 1.120 ;
  LAYER metal1 ;
  RECT 2847.720 0.000 2848.840 1.120 ;
 END
END DIA100
PIN DOA100
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2834.080 0.000 2835.200 1.120 ;
  LAYER metal4 ;
  RECT 2834.080 0.000 2835.200 1.120 ;
  LAYER metal3 ;
  RECT 2834.080 0.000 2835.200 1.120 ;
  LAYER metal2 ;
  RECT 2834.080 0.000 2835.200 1.120 ;
  LAYER metal1 ;
  RECT 2834.080 0.000 2835.200 1.120 ;
 END
END DOA100
PIN DIA99
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2820.440 0.000 2821.560 1.120 ;
  LAYER metal4 ;
  RECT 2820.440 0.000 2821.560 1.120 ;
  LAYER metal3 ;
  RECT 2820.440 0.000 2821.560 1.120 ;
  LAYER metal2 ;
  RECT 2820.440 0.000 2821.560 1.120 ;
  LAYER metal1 ;
  RECT 2820.440 0.000 2821.560 1.120 ;
 END
END DIA99
PIN DOA99
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2807.420 0.000 2808.540 1.120 ;
  LAYER metal4 ;
  RECT 2807.420 0.000 2808.540 1.120 ;
  LAYER metal3 ;
  RECT 2807.420 0.000 2808.540 1.120 ;
  LAYER metal2 ;
  RECT 2807.420 0.000 2808.540 1.120 ;
  LAYER metal1 ;
  RECT 2807.420 0.000 2808.540 1.120 ;
 END
END DOA99
PIN DIA98
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2793.780 0.000 2794.900 1.120 ;
  LAYER metal4 ;
  RECT 2793.780 0.000 2794.900 1.120 ;
  LAYER metal3 ;
  RECT 2793.780 0.000 2794.900 1.120 ;
  LAYER metal2 ;
  RECT 2793.780 0.000 2794.900 1.120 ;
  LAYER metal1 ;
  RECT 2793.780 0.000 2794.900 1.120 ;
 END
END DIA98
PIN DOA98
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2780.140 0.000 2781.260 1.120 ;
  LAYER metal4 ;
  RECT 2780.140 0.000 2781.260 1.120 ;
  LAYER metal3 ;
  RECT 2780.140 0.000 2781.260 1.120 ;
  LAYER metal2 ;
  RECT 2780.140 0.000 2781.260 1.120 ;
  LAYER metal1 ;
  RECT 2780.140 0.000 2781.260 1.120 ;
 END
END DOA98
PIN DIA97
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2767.120 0.000 2768.240 1.120 ;
  LAYER metal4 ;
  RECT 2767.120 0.000 2768.240 1.120 ;
  LAYER metal3 ;
  RECT 2767.120 0.000 2768.240 1.120 ;
  LAYER metal2 ;
  RECT 2767.120 0.000 2768.240 1.120 ;
  LAYER metal1 ;
  RECT 2767.120 0.000 2768.240 1.120 ;
 END
END DIA97
PIN DOA97
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2753.480 0.000 2754.600 1.120 ;
  LAYER metal4 ;
  RECT 2753.480 0.000 2754.600 1.120 ;
  LAYER metal3 ;
  RECT 2753.480 0.000 2754.600 1.120 ;
  LAYER metal2 ;
  RECT 2753.480 0.000 2754.600 1.120 ;
  LAYER metal1 ;
  RECT 2753.480 0.000 2754.600 1.120 ;
 END
END DOA97
PIN DIA96
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2739.840 0.000 2740.960 1.120 ;
  LAYER metal4 ;
  RECT 2739.840 0.000 2740.960 1.120 ;
  LAYER metal3 ;
  RECT 2739.840 0.000 2740.960 1.120 ;
  LAYER metal2 ;
  RECT 2739.840 0.000 2740.960 1.120 ;
  LAYER metal1 ;
  RECT 2739.840 0.000 2740.960 1.120 ;
 END
END DIA96
PIN DOA96
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2726.200 0.000 2727.320 1.120 ;
  LAYER metal4 ;
  RECT 2726.200 0.000 2727.320 1.120 ;
  LAYER metal3 ;
  RECT 2726.200 0.000 2727.320 1.120 ;
  LAYER metal2 ;
  RECT 2726.200 0.000 2727.320 1.120 ;
  LAYER metal1 ;
  RECT 2726.200 0.000 2727.320 1.120 ;
 END
END DOA96
PIN DIA95
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2713.180 0.000 2714.300 1.120 ;
  LAYER metal4 ;
  RECT 2713.180 0.000 2714.300 1.120 ;
  LAYER metal3 ;
  RECT 2713.180 0.000 2714.300 1.120 ;
  LAYER metal2 ;
  RECT 2713.180 0.000 2714.300 1.120 ;
  LAYER metal1 ;
  RECT 2713.180 0.000 2714.300 1.120 ;
 END
END DIA95
PIN DOA95
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2699.540 0.000 2700.660 1.120 ;
  LAYER metal4 ;
  RECT 2699.540 0.000 2700.660 1.120 ;
  LAYER metal3 ;
  RECT 2699.540 0.000 2700.660 1.120 ;
  LAYER metal2 ;
  RECT 2699.540 0.000 2700.660 1.120 ;
  LAYER metal1 ;
  RECT 2699.540 0.000 2700.660 1.120 ;
 END
END DOA95
PIN DIA94
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2685.900 0.000 2687.020 1.120 ;
  LAYER metal4 ;
  RECT 2685.900 0.000 2687.020 1.120 ;
  LAYER metal3 ;
  RECT 2685.900 0.000 2687.020 1.120 ;
  LAYER metal2 ;
  RECT 2685.900 0.000 2687.020 1.120 ;
  LAYER metal1 ;
  RECT 2685.900 0.000 2687.020 1.120 ;
 END
END DIA94
PIN DOA94
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2672.880 0.000 2674.000 1.120 ;
  LAYER metal4 ;
  RECT 2672.880 0.000 2674.000 1.120 ;
  LAYER metal3 ;
  RECT 2672.880 0.000 2674.000 1.120 ;
  LAYER metal2 ;
  RECT 2672.880 0.000 2674.000 1.120 ;
  LAYER metal1 ;
  RECT 2672.880 0.000 2674.000 1.120 ;
 END
END DOA94
PIN DIA93
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2659.240 0.000 2660.360 1.120 ;
  LAYER metal4 ;
  RECT 2659.240 0.000 2660.360 1.120 ;
  LAYER metal3 ;
  RECT 2659.240 0.000 2660.360 1.120 ;
  LAYER metal2 ;
  RECT 2659.240 0.000 2660.360 1.120 ;
  LAYER metal1 ;
  RECT 2659.240 0.000 2660.360 1.120 ;
 END
END DIA93
PIN DOA93
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2645.600 0.000 2646.720 1.120 ;
  LAYER metal4 ;
  RECT 2645.600 0.000 2646.720 1.120 ;
  LAYER metal3 ;
  RECT 2645.600 0.000 2646.720 1.120 ;
  LAYER metal2 ;
  RECT 2645.600 0.000 2646.720 1.120 ;
  LAYER metal1 ;
  RECT 2645.600 0.000 2646.720 1.120 ;
 END
END DOA93
PIN DIA92
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2632.580 0.000 2633.700 1.120 ;
  LAYER metal4 ;
  RECT 2632.580 0.000 2633.700 1.120 ;
  LAYER metal3 ;
  RECT 2632.580 0.000 2633.700 1.120 ;
  LAYER metal2 ;
  RECT 2632.580 0.000 2633.700 1.120 ;
  LAYER metal1 ;
  RECT 2632.580 0.000 2633.700 1.120 ;
 END
END DIA92
PIN DOA92
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2618.940 0.000 2620.060 1.120 ;
  LAYER metal4 ;
  RECT 2618.940 0.000 2620.060 1.120 ;
  LAYER metal3 ;
  RECT 2618.940 0.000 2620.060 1.120 ;
  LAYER metal2 ;
  RECT 2618.940 0.000 2620.060 1.120 ;
  LAYER metal1 ;
  RECT 2618.940 0.000 2620.060 1.120 ;
 END
END DOA92
PIN DIA91
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2605.300 0.000 2606.420 1.120 ;
  LAYER metal4 ;
  RECT 2605.300 0.000 2606.420 1.120 ;
  LAYER metal3 ;
  RECT 2605.300 0.000 2606.420 1.120 ;
  LAYER metal2 ;
  RECT 2605.300 0.000 2606.420 1.120 ;
  LAYER metal1 ;
  RECT 2605.300 0.000 2606.420 1.120 ;
 END
END DIA91
PIN DOA91
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2592.280 0.000 2593.400 1.120 ;
  LAYER metal4 ;
  RECT 2592.280 0.000 2593.400 1.120 ;
  LAYER metal3 ;
  RECT 2592.280 0.000 2593.400 1.120 ;
  LAYER metal2 ;
  RECT 2592.280 0.000 2593.400 1.120 ;
  LAYER metal1 ;
  RECT 2592.280 0.000 2593.400 1.120 ;
 END
END DOA91
PIN DIA90
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2578.640 0.000 2579.760 1.120 ;
  LAYER metal4 ;
  RECT 2578.640 0.000 2579.760 1.120 ;
  LAYER metal3 ;
  RECT 2578.640 0.000 2579.760 1.120 ;
  LAYER metal2 ;
  RECT 2578.640 0.000 2579.760 1.120 ;
  LAYER metal1 ;
  RECT 2578.640 0.000 2579.760 1.120 ;
 END
END DIA90
PIN DOA90
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2565.000 0.000 2566.120 1.120 ;
  LAYER metal4 ;
  RECT 2565.000 0.000 2566.120 1.120 ;
  LAYER metal3 ;
  RECT 2565.000 0.000 2566.120 1.120 ;
  LAYER metal2 ;
  RECT 2565.000 0.000 2566.120 1.120 ;
  LAYER metal1 ;
  RECT 2565.000 0.000 2566.120 1.120 ;
 END
END DOA90
PIN DIA89
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2551.980 0.000 2553.100 1.120 ;
  LAYER metal4 ;
  RECT 2551.980 0.000 2553.100 1.120 ;
  LAYER metal3 ;
  RECT 2551.980 0.000 2553.100 1.120 ;
  LAYER metal2 ;
  RECT 2551.980 0.000 2553.100 1.120 ;
  LAYER metal1 ;
  RECT 2551.980 0.000 2553.100 1.120 ;
 END
END DIA89
PIN DOA89
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2538.340 0.000 2539.460 1.120 ;
  LAYER metal4 ;
  RECT 2538.340 0.000 2539.460 1.120 ;
  LAYER metal3 ;
  RECT 2538.340 0.000 2539.460 1.120 ;
  LAYER metal2 ;
  RECT 2538.340 0.000 2539.460 1.120 ;
  LAYER metal1 ;
  RECT 2538.340 0.000 2539.460 1.120 ;
 END
END DOA89
PIN DIA88
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2524.700 0.000 2525.820 1.120 ;
  LAYER metal4 ;
  RECT 2524.700 0.000 2525.820 1.120 ;
  LAYER metal3 ;
  RECT 2524.700 0.000 2525.820 1.120 ;
  LAYER metal2 ;
  RECT 2524.700 0.000 2525.820 1.120 ;
  LAYER metal1 ;
  RECT 2524.700 0.000 2525.820 1.120 ;
 END
END DIA88
PIN DOA88
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2511.680 0.000 2512.800 1.120 ;
  LAYER metal4 ;
  RECT 2511.680 0.000 2512.800 1.120 ;
  LAYER metal3 ;
  RECT 2511.680 0.000 2512.800 1.120 ;
  LAYER metal2 ;
  RECT 2511.680 0.000 2512.800 1.120 ;
  LAYER metal1 ;
  RECT 2511.680 0.000 2512.800 1.120 ;
 END
END DOA88
PIN DIA87
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2498.040 0.000 2499.160 1.120 ;
  LAYER metal4 ;
  RECT 2498.040 0.000 2499.160 1.120 ;
  LAYER metal3 ;
  RECT 2498.040 0.000 2499.160 1.120 ;
  LAYER metal2 ;
  RECT 2498.040 0.000 2499.160 1.120 ;
  LAYER metal1 ;
  RECT 2498.040 0.000 2499.160 1.120 ;
 END
END DIA87
PIN DOA87
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2484.400 0.000 2485.520 1.120 ;
  LAYER metal4 ;
  RECT 2484.400 0.000 2485.520 1.120 ;
  LAYER metal3 ;
  RECT 2484.400 0.000 2485.520 1.120 ;
  LAYER metal2 ;
  RECT 2484.400 0.000 2485.520 1.120 ;
  LAYER metal1 ;
  RECT 2484.400 0.000 2485.520 1.120 ;
 END
END DOA87
PIN DIA86
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2471.380 0.000 2472.500 1.120 ;
  LAYER metal4 ;
  RECT 2471.380 0.000 2472.500 1.120 ;
  LAYER metal3 ;
  RECT 2471.380 0.000 2472.500 1.120 ;
  LAYER metal2 ;
  RECT 2471.380 0.000 2472.500 1.120 ;
  LAYER metal1 ;
  RECT 2471.380 0.000 2472.500 1.120 ;
 END
END DIA86
PIN DOA86
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2457.740 0.000 2458.860 1.120 ;
  LAYER metal4 ;
  RECT 2457.740 0.000 2458.860 1.120 ;
  LAYER metal3 ;
  RECT 2457.740 0.000 2458.860 1.120 ;
  LAYER metal2 ;
  RECT 2457.740 0.000 2458.860 1.120 ;
  LAYER metal1 ;
  RECT 2457.740 0.000 2458.860 1.120 ;
 END
END DOA86
PIN DIA85
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2444.100 0.000 2445.220 1.120 ;
  LAYER metal4 ;
  RECT 2444.100 0.000 2445.220 1.120 ;
  LAYER metal3 ;
  RECT 2444.100 0.000 2445.220 1.120 ;
  LAYER metal2 ;
  RECT 2444.100 0.000 2445.220 1.120 ;
  LAYER metal1 ;
  RECT 2444.100 0.000 2445.220 1.120 ;
 END
END DIA85
PIN DOA85
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2431.080 0.000 2432.200 1.120 ;
  LAYER metal4 ;
  RECT 2431.080 0.000 2432.200 1.120 ;
  LAYER metal3 ;
  RECT 2431.080 0.000 2432.200 1.120 ;
  LAYER metal2 ;
  RECT 2431.080 0.000 2432.200 1.120 ;
  LAYER metal1 ;
  RECT 2431.080 0.000 2432.200 1.120 ;
 END
END DOA85
PIN DIA84
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2417.440 0.000 2418.560 1.120 ;
  LAYER metal4 ;
  RECT 2417.440 0.000 2418.560 1.120 ;
  LAYER metal3 ;
  RECT 2417.440 0.000 2418.560 1.120 ;
  LAYER metal2 ;
  RECT 2417.440 0.000 2418.560 1.120 ;
  LAYER metal1 ;
  RECT 2417.440 0.000 2418.560 1.120 ;
 END
END DIA84
PIN DOA84
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2403.800 0.000 2404.920 1.120 ;
  LAYER metal4 ;
  RECT 2403.800 0.000 2404.920 1.120 ;
  LAYER metal3 ;
  RECT 2403.800 0.000 2404.920 1.120 ;
  LAYER metal2 ;
  RECT 2403.800 0.000 2404.920 1.120 ;
  LAYER metal1 ;
  RECT 2403.800 0.000 2404.920 1.120 ;
 END
END DOA84
PIN DIA83
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2390.780 0.000 2391.900 1.120 ;
  LAYER metal4 ;
  RECT 2390.780 0.000 2391.900 1.120 ;
  LAYER metal3 ;
  RECT 2390.780 0.000 2391.900 1.120 ;
  LAYER metal2 ;
  RECT 2390.780 0.000 2391.900 1.120 ;
  LAYER metal1 ;
  RECT 2390.780 0.000 2391.900 1.120 ;
 END
END DIA83
PIN DOA83
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2377.140 0.000 2378.260 1.120 ;
  LAYER metal4 ;
  RECT 2377.140 0.000 2378.260 1.120 ;
  LAYER metal3 ;
  RECT 2377.140 0.000 2378.260 1.120 ;
  LAYER metal2 ;
  RECT 2377.140 0.000 2378.260 1.120 ;
  LAYER metal1 ;
  RECT 2377.140 0.000 2378.260 1.120 ;
 END
END DOA83
PIN DIA82
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2363.500 0.000 2364.620 1.120 ;
  LAYER metal4 ;
  RECT 2363.500 0.000 2364.620 1.120 ;
  LAYER metal3 ;
  RECT 2363.500 0.000 2364.620 1.120 ;
  LAYER metal2 ;
  RECT 2363.500 0.000 2364.620 1.120 ;
  LAYER metal1 ;
  RECT 2363.500 0.000 2364.620 1.120 ;
 END
END DIA82
PIN DOA82
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2350.480 0.000 2351.600 1.120 ;
  LAYER metal4 ;
  RECT 2350.480 0.000 2351.600 1.120 ;
  LAYER metal3 ;
  RECT 2350.480 0.000 2351.600 1.120 ;
  LAYER metal2 ;
  RECT 2350.480 0.000 2351.600 1.120 ;
  LAYER metal1 ;
  RECT 2350.480 0.000 2351.600 1.120 ;
 END
END DOA82
PIN DIA81
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2336.840 0.000 2337.960 1.120 ;
  LAYER metal4 ;
  RECT 2336.840 0.000 2337.960 1.120 ;
  LAYER metal3 ;
  RECT 2336.840 0.000 2337.960 1.120 ;
  LAYER metal2 ;
  RECT 2336.840 0.000 2337.960 1.120 ;
  LAYER metal1 ;
  RECT 2336.840 0.000 2337.960 1.120 ;
 END
END DIA81
PIN DOA81
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2323.200 0.000 2324.320 1.120 ;
  LAYER metal4 ;
  RECT 2323.200 0.000 2324.320 1.120 ;
  LAYER metal3 ;
  RECT 2323.200 0.000 2324.320 1.120 ;
  LAYER metal2 ;
  RECT 2323.200 0.000 2324.320 1.120 ;
  LAYER metal1 ;
  RECT 2323.200 0.000 2324.320 1.120 ;
 END
END DOA81
PIN DIA80
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2309.560 0.000 2310.680 1.120 ;
  LAYER metal4 ;
  RECT 2309.560 0.000 2310.680 1.120 ;
  LAYER metal3 ;
  RECT 2309.560 0.000 2310.680 1.120 ;
  LAYER metal2 ;
  RECT 2309.560 0.000 2310.680 1.120 ;
  LAYER metal1 ;
  RECT 2309.560 0.000 2310.680 1.120 ;
 END
END DIA80
PIN DOA80
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2296.540 0.000 2297.660 1.120 ;
  LAYER metal4 ;
  RECT 2296.540 0.000 2297.660 1.120 ;
  LAYER metal3 ;
  RECT 2296.540 0.000 2297.660 1.120 ;
  LAYER metal2 ;
  RECT 2296.540 0.000 2297.660 1.120 ;
  LAYER metal1 ;
  RECT 2296.540 0.000 2297.660 1.120 ;
 END
END DOA80
PIN DIA79
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2282.900 0.000 2284.020 1.120 ;
  LAYER metal4 ;
  RECT 2282.900 0.000 2284.020 1.120 ;
  LAYER metal3 ;
  RECT 2282.900 0.000 2284.020 1.120 ;
  LAYER metal2 ;
  RECT 2282.900 0.000 2284.020 1.120 ;
  LAYER metal1 ;
  RECT 2282.900 0.000 2284.020 1.120 ;
 END
END DIA79
PIN DOA79
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2269.260 0.000 2270.380 1.120 ;
  LAYER metal4 ;
  RECT 2269.260 0.000 2270.380 1.120 ;
  LAYER metal3 ;
  RECT 2269.260 0.000 2270.380 1.120 ;
  LAYER metal2 ;
  RECT 2269.260 0.000 2270.380 1.120 ;
  LAYER metal1 ;
  RECT 2269.260 0.000 2270.380 1.120 ;
 END
END DOA79
PIN DIA78
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2256.240 0.000 2257.360 1.120 ;
  LAYER metal4 ;
  RECT 2256.240 0.000 2257.360 1.120 ;
  LAYER metal3 ;
  RECT 2256.240 0.000 2257.360 1.120 ;
  LAYER metal2 ;
  RECT 2256.240 0.000 2257.360 1.120 ;
  LAYER metal1 ;
  RECT 2256.240 0.000 2257.360 1.120 ;
 END
END DIA78
PIN DOA78
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2242.600 0.000 2243.720 1.120 ;
  LAYER metal4 ;
  RECT 2242.600 0.000 2243.720 1.120 ;
  LAYER metal3 ;
  RECT 2242.600 0.000 2243.720 1.120 ;
  LAYER metal2 ;
  RECT 2242.600 0.000 2243.720 1.120 ;
  LAYER metal1 ;
  RECT 2242.600 0.000 2243.720 1.120 ;
 END
END DOA78
PIN DIA77
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2228.960 0.000 2230.080 1.120 ;
  LAYER metal4 ;
  RECT 2228.960 0.000 2230.080 1.120 ;
  LAYER metal3 ;
  RECT 2228.960 0.000 2230.080 1.120 ;
  LAYER metal2 ;
  RECT 2228.960 0.000 2230.080 1.120 ;
  LAYER metal1 ;
  RECT 2228.960 0.000 2230.080 1.120 ;
 END
END DIA77
PIN DOA77
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2215.940 0.000 2217.060 1.120 ;
  LAYER metal4 ;
  RECT 2215.940 0.000 2217.060 1.120 ;
  LAYER metal3 ;
  RECT 2215.940 0.000 2217.060 1.120 ;
  LAYER metal2 ;
  RECT 2215.940 0.000 2217.060 1.120 ;
  LAYER metal1 ;
  RECT 2215.940 0.000 2217.060 1.120 ;
 END
END DOA77
PIN DIA76
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2202.300 0.000 2203.420 1.120 ;
  LAYER metal4 ;
  RECT 2202.300 0.000 2203.420 1.120 ;
  LAYER metal3 ;
  RECT 2202.300 0.000 2203.420 1.120 ;
  LAYER metal2 ;
  RECT 2202.300 0.000 2203.420 1.120 ;
  LAYER metal1 ;
  RECT 2202.300 0.000 2203.420 1.120 ;
 END
END DIA76
PIN DOA76
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2188.660 0.000 2189.780 1.120 ;
  LAYER metal4 ;
  RECT 2188.660 0.000 2189.780 1.120 ;
  LAYER metal3 ;
  RECT 2188.660 0.000 2189.780 1.120 ;
  LAYER metal2 ;
  RECT 2188.660 0.000 2189.780 1.120 ;
  LAYER metal1 ;
  RECT 2188.660 0.000 2189.780 1.120 ;
 END
END DOA76
PIN DIA75
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2175.640 0.000 2176.760 1.120 ;
  LAYER metal4 ;
  RECT 2175.640 0.000 2176.760 1.120 ;
  LAYER metal3 ;
  RECT 2175.640 0.000 2176.760 1.120 ;
  LAYER metal2 ;
  RECT 2175.640 0.000 2176.760 1.120 ;
  LAYER metal1 ;
  RECT 2175.640 0.000 2176.760 1.120 ;
 END
END DIA75
PIN DOA75
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2162.000 0.000 2163.120 1.120 ;
  LAYER metal4 ;
  RECT 2162.000 0.000 2163.120 1.120 ;
  LAYER metal3 ;
  RECT 2162.000 0.000 2163.120 1.120 ;
  LAYER metal2 ;
  RECT 2162.000 0.000 2163.120 1.120 ;
  LAYER metal1 ;
  RECT 2162.000 0.000 2163.120 1.120 ;
 END
END DOA75
PIN DIA74
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2148.360 0.000 2149.480 1.120 ;
  LAYER metal4 ;
  RECT 2148.360 0.000 2149.480 1.120 ;
  LAYER metal3 ;
  RECT 2148.360 0.000 2149.480 1.120 ;
  LAYER metal2 ;
  RECT 2148.360 0.000 2149.480 1.120 ;
  LAYER metal1 ;
  RECT 2148.360 0.000 2149.480 1.120 ;
 END
END DIA74
PIN DOA74
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2135.340 0.000 2136.460 1.120 ;
  LAYER metal4 ;
  RECT 2135.340 0.000 2136.460 1.120 ;
  LAYER metal3 ;
  RECT 2135.340 0.000 2136.460 1.120 ;
  LAYER metal2 ;
  RECT 2135.340 0.000 2136.460 1.120 ;
  LAYER metal1 ;
  RECT 2135.340 0.000 2136.460 1.120 ;
 END
END DOA74
PIN DIA73
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2121.700 0.000 2122.820 1.120 ;
  LAYER metal4 ;
  RECT 2121.700 0.000 2122.820 1.120 ;
  LAYER metal3 ;
  RECT 2121.700 0.000 2122.820 1.120 ;
  LAYER metal2 ;
  RECT 2121.700 0.000 2122.820 1.120 ;
  LAYER metal1 ;
  RECT 2121.700 0.000 2122.820 1.120 ;
 END
END DIA73
PIN DOA73
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2108.060 0.000 2109.180 1.120 ;
  LAYER metal4 ;
  RECT 2108.060 0.000 2109.180 1.120 ;
  LAYER metal3 ;
  RECT 2108.060 0.000 2109.180 1.120 ;
  LAYER metal2 ;
  RECT 2108.060 0.000 2109.180 1.120 ;
  LAYER metal1 ;
  RECT 2108.060 0.000 2109.180 1.120 ;
 END
END DOA73
PIN DIA72
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2095.040 0.000 2096.160 1.120 ;
  LAYER metal4 ;
  RECT 2095.040 0.000 2096.160 1.120 ;
  LAYER metal3 ;
  RECT 2095.040 0.000 2096.160 1.120 ;
  LAYER metal2 ;
  RECT 2095.040 0.000 2096.160 1.120 ;
  LAYER metal1 ;
  RECT 2095.040 0.000 2096.160 1.120 ;
 END
END DIA72
PIN DOA72
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2081.400 0.000 2082.520 1.120 ;
  LAYER metal4 ;
  RECT 2081.400 0.000 2082.520 1.120 ;
  LAYER metal3 ;
  RECT 2081.400 0.000 2082.520 1.120 ;
  LAYER metal2 ;
  RECT 2081.400 0.000 2082.520 1.120 ;
  LAYER metal1 ;
  RECT 2081.400 0.000 2082.520 1.120 ;
 END
END DOA72
PIN DIA71
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2067.760 0.000 2068.880 1.120 ;
  LAYER metal4 ;
  RECT 2067.760 0.000 2068.880 1.120 ;
  LAYER metal3 ;
  RECT 2067.760 0.000 2068.880 1.120 ;
  LAYER metal2 ;
  RECT 2067.760 0.000 2068.880 1.120 ;
  LAYER metal1 ;
  RECT 2067.760 0.000 2068.880 1.120 ;
 END
END DIA71
PIN DOA71
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2054.740 0.000 2055.860 1.120 ;
  LAYER metal4 ;
  RECT 2054.740 0.000 2055.860 1.120 ;
  LAYER metal3 ;
  RECT 2054.740 0.000 2055.860 1.120 ;
  LAYER metal2 ;
  RECT 2054.740 0.000 2055.860 1.120 ;
  LAYER metal1 ;
  RECT 2054.740 0.000 2055.860 1.120 ;
 END
END DOA71
PIN DIA70
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2041.100 0.000 2042.220 1.120 ;
  LAYER metal4 ;
  RECT 2041.100 0.000 2042.220 1.120 ;
  LAYER metal3 ;
  RECT 2041.100 0.000 2042.220 1.120 ;
  LAYER metal2 ;
  RECT 2041.100 0.000 2042.220 1.120 ;
  LAYER metal1 ;
  RECT 2041.100 0.000 2042.220 1.120 ;
 END
END DIA70
PIN DOA70
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2027.460 0.000 2028.580 1.120 ;
  LAYER metal4 ;
  RECT 2027.460 0.000 2028.580 1.120 ;
  LAYER metal3 ;
  RECT 2027.460 0.000 2028.580 1.120 ;
  LAYER metal2 ;
  RECT 2027.460 0.000 2028.580 1.120 ;
  LAYER metal1 ;
  RECT 2027.460 0.000 2028.580 1.120 ;
 END
END DOA70
PIN DIA69
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2014.440 0.000 2015.560 1.120 ;
  LAYER metal4 ;
  RECT 2014.440 0.000 2015.560 1.120 ;
  LAYER metal3 ;
  RECT 2014.440 0.000 2015.560 1.120 ;
  LAYER metal2 ;
  RECT 2014.440 0.000 2015.560 1.120 ;
  LAYER metal1 ;
  RECT 2014.440 0.000 2015.560 1.120 ;
 END
END DIA69
PIN DOA69
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2000.800 0.000 2001.920 1.120 ;
  LAYER metal4 ;
  RECT 2000.800 0.000 2001.920 1.120 ;
  LAYER metal3 ;
  RECT 2000.800 0.000 2001.920 1.120 ;
  LAYER metal2 ;
  RECT 2000.800 0.000 2001.920 1.120 ;
  LAYER metal1 ;
  RECT 2000.800 0.000 2001.920 1.120 ;
 END
END DOA69
PIN DIA68
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1987.160 0.000 1988.280 1.120 ;
  LAYER metal4 ;
  RECT 1987.160 0.000 1988.280 1.120 ;
  LAYER metal3 ;
  RECT 1987.160 0.000 1988.280 1.120 ;
  LAYER metal2 ;
  RECT 1987.160 0.000 1988.280 1.120 ;
  LAYER metal1 ;
  RECT 1987.160 0.000 1988.280 1.120 ;
 END
END DIA68
PIN DOA68
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1974.140 0.000 1975.260 1.120 ;
  LAYER metal4 ;
  RECT 1974.140 0.000 1975.260 1.120 ;
  LAYER metal3 ;
  RECT 1974.140 0.000 1975.260 1.120 ;
  LAYER metal2 ;
  RECT 1974.140 0.000 1975.260 1.120 ;
  LAYER metal1 ;
  RECT 1974.140 0.000 1975.260 1.120 ;
 END
END DOA68
PIN DIA67
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1960.500 0.000 1961.620 1.120 ;
  LAYER metal4 ;
  RECT 1960.500 0.000 1961.620 1.120 ;
  LAYER metal3 ;
  RECT 1960.500 0.000 1961.620 1.120 ;
  LAYER metal2 ;
  RECT 1960.500 0.000 1961.620 1.120 ;
  LAYER metal1 ;
  RECT 1960.500 0.000 1961.620 1.120 ;
 END
END DIA67
PIN DOA67
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1946.860 0.000 1947.980 1.120 ;
  LAYER metal4 ;
  RECT 1946.860 0.000 1947.980 1.120 ;
  LAYER metal3 ;
  RECT 1946.860 0.000 1947.980 1.120 ;
  LAYER metal2 ;
  RECT 1946.860 0.000 1947.980 1.120 ;
  LAYER metal1 ;
  RECT 1946.860 0.000 1947.980 1.120 ;
 END
END DOA67
PIN DIA66
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1933.840 0.000 1934.960 1.120 ;
  LAYER metal4 ;
  RECT 1933.840 0.000 1934.960 1.120 ;
  LAYER metal3 ;
  RECT 1933.840 0.000 1934.960 1.120 ;
  LAYER metal2 ;
  RECT 1933.840 0.000 1934.960 1.120 ;
  LAYER metal1 ;
  RECT 1933.840 0.000 1934.960 1.120 ;
 END
END DIA66
PIN DOA66
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1920.200 0.000 1921.320 1.120 ;
  LAYER metal4 ;
  RECT 1920.200 0.000 1921.320 1.120 ;
  LAYER metal3 ;
  RECT 1920.200 0.000 1921.320 1.120 ;
  LAYER metal2 ;
  RECT 1920.200 0.000 1921.320 1.120 ;
  LAYER metal1 ;
  RECT 1920.200 0.000 1921.320 1.120 ;
 END
END DOA66
PIN DIA65
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1906.560 0.000 1907.680 1.120 ;
  LAYER metal4 ;
  RECT 1906.560 0.000 1907.680 1.120 ;
  LAYER metal3 ;
  RECT 1906.560 0.000 1907.680 1.120 ;
  LAYER metal2 ;
  RECT 1906.560 0.000 1907.680 1.120 ;
  LAYER metal1 ;
  RECT 1906.560 0.000 1907.680 1.120 ;
 END
END DIA65
PIN DOA65
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1892.920 0.000 1894.040 1.120 ;
  LAYER metal4 ;
  RECT 1892.920 0.000 1894.040 1.120 ;
  LAYER metal3 ;
  RECT 1892.920 0.000 1894.040 1.120 ;
  LAYER metal2 ;
  RECT 1892.920 0.000 1894.040 1.120 ;
  LAYER metal1 ;
  RECT 1892.920 0.000 1894.040 1.120 ;
 END
END DOA65
PIN DIA64
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1879.900 0.000 1881.020 1.120 ;
  LAYER metal4 ;
  RECT 1879.900 0.000 1881.020 1.120 ;
  LAYER metal3 ;
  RECT 1879.900 0.000 1881.020 1.120 ;
  LAYER metal2 ;
  RECT 1879.900 0.000 1881.020 1.120 ;
  LAYER metal1 ;
  RECT 1879.900 0.000 1881.020 1.120 ;
 END
END DIA64
PIN DOA64
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1866.260 0.000 1867.380 1.120 ;
  LAYER metal4 ;
  RECT 1866.260 0.000 1867.380 1.120 ;
  LAYER metal3 ;
  RECT 1866.260 0.000 1867.380 1.120 ;
  LAYER metal2 ;
  RECT 1866.260 0.000 1867.380 1.120 ;
  LAYER metal1 ;
  RECT 1866.260 0.000 1867.380 1.120 ;
 END
END DOA64
PIN OEA
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1839.600 0.000 1840.720 1.120 ;
  LAYER metal4 ;
  RECT 1839.600 0.000 1840.720 1.120 ;
  LAYER metal3 ;
  RECT 1839.600 0.000 1840.720 1.120 ;
  LAYER metal2 ;
  RECT 1839.600 0.000 1840.720 1.120 ;
  LAYER metal1 ;
  RECT 1839.600 0.000 1840.720 1.120 ;
 END
END OEA
PIN CKA
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1826.580 0.000 1827.700 1.120 ;
  LAYER metal4 ;
  RECT 1826.580 0.000 1827.700 1.120 ;
  LAYER metal3 ;
  RECT 1826.580 0.000 1827.700 1.120 ;
  LAYER metal2 ;
  RECT 1826.580 0.000 1827.700 1.120 ;
  LAYER metal1 ;
  RECT 1826.580 0.000 1827.700 1.120 ;
 END
END CKA
PIN CSA
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1824.720 0.000 1825.840 1.120 ;
  LAYER metal4 ;
  RECT 1824.720 0.000 1825.840 1.120 ;
  LAYER metal3 ;
  RECT 1824.720 0.000 1825.840 1.120 ;
  LAYER metal2 ;
  RECT 1824.720 0.000 1825.840 1.120 ;
  LAYER metal1 ;
  RECT 1824.720 0.000 1825.840 1.120 ;
 END
END CSA
PIN WEAN
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1821.620 0.000 1822.740 1.120 ;
  LAYER metal4 ;
  RECT 1821.620 0.000 1822.740 1.120 ;
  LAYER metal3 ;
  RECT 1821.620 0.000 1822.740 1.120 ;
  LAYER metal2 ;
  RECT 1821.620 0.000 1822.740 1.120 ;
  LAYER metal1 ;
  RECT 1821.620 0.000 1822.740 1.120 ;
 END
END WEAN
PIN A2
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1817.900 0.000 1819.020 1.120 ;
  LAYER metal4 ;
  RECT 1817.900 0.000 1819.020 1.120 ;
  LAYER metal3 ;
  RECT 1817.900 0.000 1819.020 1.120 ;
  LAYER metal2 ;
  RECT 1817.900 0.000 1819.020 1.120 ;
  LAYER metal1 ;
  RECT 1817.900 0.000 1819.020 1.120 ;
 END
END A2
PIN A1
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1812.940 0.000 1814.060 1.120 ;
  LAYER metal4 ;
  RECT 1812.940 0.000 1814.060 1.120 ;
  LAYER metal3 ;
  RECT 1812.940 0.000 1814.060 1.120 ;
  LAYER metal2 ;
  RECT 1812.940 0.000 1814.060 1.120 ;
  LAYER metal1 ;
  RECT 1812.940 0.000 1814.060 1.120 ;
 END
END A1
PIN A0
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1810.460 0.000 1811.580 1.120 ;
  LAYER metal4 ;
  RECT 1810.460 0.000 1811.580 1.120 ;
  LAYER metal3 ;
  RECT 1810.460 0.000 1811.580 1.120 ;
  LAYER metal2 ;
  RECT 1810.460 0.000 1811.580 1.120 ;
  LAYER metal1 ;
  RECT 1810.460 0.000 1811.580 1.120 ;
 END
END A0
PIN A5
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1801.780 0.000 1802.900 1.120 ;
  LAYER metal4 ;
  RECT 1801.780 0.000 1802.900 1.120 ;
  LAYER metal3 ;
  RECT 1801.780 0.000 1802.900 1.120 ;
  LAYER metal2 ;
  RECT 1801.780 0.000 1802.900 1.120 ;
  LAYER metal1 ;
  RECT 1801.780 0.000 1802.900 1.120 ;
 END
END A5
PIN A4
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1796.200 0.000 1797.320 1.120 ;
  LAYER metal4 ;
  RECT 1796.200 0.000 1797.320 1.120 ;
  LAYER metal3 ;
  RECT 1796.200 0.000 1797.320 1.120 ;
  LAYER metal2 ;
  RECT 1796.200 0.000 1797.320 1.120 ;
  LAYER metal1 ;
  RECT 1796.200 0.000 1797.320 1.120 ;
 END
END A4
PIN A3
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1790.620 0.000 1791.740 1.120 ;
  LAYER metal4 ;
  RECT 1790.620 0.000 1791.740 1.120 ;
  LAYER metal3 ;
  RECT 1790.620 0.000 1791.740 1.120 ;
  LAYER metal2 ;
  RECT 1790.620 0.000 1791.740 1.120 ;
  LAYER metal1 ;
  RECT 1790.620 0.000 1791.740 1.120 ;
 END
END A3
PIN A8
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1777.600 0.000 1778.720 1.120 ;
  LAYER metal4 ;
  RECT 1777.600 0.000 1778.720 1.120 ;
  LAYER metal3 ;
  RECT 1777.600 0.000 1778.720 1.120 ;
  LAYER metal2 ;
  RECT 1777.600 0.000 1778.720 1.120 ;
  LAYER metal1 ;
  RECT 1777.600 0.000 1778.720 1.120 ;
 END
END A8
PIN A7
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1772.020 0.000 1773.140 1.120 ;
  LAYER metal4 ;
  RECT 1772.020 0.000 1773.140 1.120 ;
  LAYER metal3 ;
  RECT 1772.020 0.000 1773.140 1.120 ;
  LAYER metal2 ;
  RECT 1772.020 0.000 1773.140 1.120 ;
  LAYER metal1 ;
  RECT 1772.020 0.000 1773.140 1.120 ;
 END
END A7
PIN A6
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1766.440 0.000 1767.560 1.120 ;
  LAYER metal4 ;
  RECT 1766.440 0.000 1767.560 1.120 ;
  LAYER metal3 ;
  RECT 1766.440 0.000 1767.560 1.120 ;
  LAYER metal2 ;
  RECT 1766.440 0.000 1767.560 1.120 ;
  LAYER metal1 ;
  RECT 1766.440 0.000 1767.560 1.120 ;
 END
END A6
PIN A9
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1741.640 0.000 1742.760 1.120 ;
  LAYER metal4 ;
  RECT 1741.640 0.000 1742.760 1.120 ;
  LAYER metal3 ;
  RECT 1741.640 0.000 1742.760 1.120 ;
  LAYER metal2 ;
  RECT 1741.640 0.000 1742.760 1.120 ;
  LAYER metal1 ;
  RECT 1741.640 0.000 1742.760 1.120 ;
 END
END A9
PIN DIA63
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1719.320 0.000 1720.440 1.120 ;
  LAYER metal4 ;
  RECT 1719.320 0.000 1720.440 1.120 ;
  LAYER metal3 ;
  RECT 1719.320 0.000 1720.440 1.120 ;
  LAYER metal2 ;
  RECT 1719.320 0.000 1720.440 1.120 ;
  LAYER metal1 ;
  RECT 1719.320 0.000 1720.440 1.120 ;
 END
END DIA63
PIN DOA63
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1706.300 0.000 1707.420 1.120 ;
  LAYER metal4 ;
  RECT 1706.300 0.000 1707.420 1.120 ;
  LAYER metal3 ;
  RECT 1706.300 0.000 1707.420 1.120 ;
  LAYER metal2 ;
  RECT 1706.300 0.000 1707.420 1.120 ;
  LAYER metal1 ;
  RECT 1706.300 0.000 1707.420 1.120 ;
 END
END DOA63
PIN DIA62
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1692.660 0.000 1693.780 1.120 ;
  LAYER metal4 ;
  RECT 1692.660 0.000 1693.780 1.120 ;
  LAYER metal3 ;
  RECT 1692.660 0.000 1693.780 1.120 ;
  LAYER metal2 ;
  RECT 1692.660 0.000 1693.780 1.120 ;
  LAYER metal1 ;
  RECT 1692.660 0.000 1693.780 1.120 ;
 END
END DIA62
PIN DOA62
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1679.020 0.000 1680.140 1.120 ;
  LAYER metal4 ;
  RECT 1679.020 0.000 1680.140 1.120 ;
  LAYER metal3 ;
  RECT 1679.020 0.000 1680.140 1.120 ;
  LAYER metal2 ;
  RECT 1679.020 0.000 1680.140 1.120 ;
  LAYER metal1 ;
  RECT 1679.020 0.000 1680.140 1.120 ;
 END
END DOA62
PIN DIA61
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1666.000 0.000 1667.120 1.120 ;
  LAYER metal4 ;
  RECT 1666.000 0.000 1667.120 1.120 ;
  LAYER metal3 ;
  RECT 1666.000 0.000 1667.120 1.120 ;
  LAYER metal2 ;
  RECT 1666.000 0.000 1667.120 1.120 ;
  LAYER metal1 ;
  RECT 1666.000 0.000 1667.120 1.120 ;
 END
END DIA61
PIN DOA61
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1652.360 0.000 1653.480 1.120 ;
  LAYER metal4 ;
  RECT 1652.360 0.000 1653.480 1.120 ;
  LAYER metal3 ;
  RECT 1652.360 0.000 1653.480 1.120 ;
  LAYER metal2 ;
  RECT 1652.360 0.000 1653.480 1.120 ;
  LAYER metal1 ;
  RECT 1652.360 0.000 1653.480 1.120 ;
 END
END DOA61
PIN DIA60
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1638.720 0.000 1639.840 1.120 ;
  LAYER metal4 ;
  RECT 1638.720 0.000 1639.840 1.120 ;
  LAYER metal3 ;
  RECT 1638.720 0.000 1639.840 1.120 ;
  LAYER metal2 ;
  RECT 1638.720 0.000 1639.840 1.120 ;
  LAYER metal1 ;
  RECT 1638.720 0.000 1639.840 1.120 ;
 END
END DIA60
PIN DOA60
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1625.700 0.000 1626.820 1.120 ;
  LAYER metal4 ;
  RECT 1625.700 0.000 1626.820 1.120 ;
  LAYER metal3 ;
  RECT 1625.700 0.000 1626.820 1.120 ;
  LAYER metal2 ;
  RECT 1625.700 0.000 1626.820 1.120 ;
  LAYER metal1 ;
  RECT 1625.700 0.000 1626.820 1.120 ;
 END
END DOA60
PIN DIA59
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1612.060 0.000 1613.180 1.120 ;
  LAYER metal4 ;
  RECT 1612.060 0.000 1613.180 1.120 ;
  LAYER metal3 ;
  RECT 1612.060 0.000 1613.180 1.120 ;
  LAYER metal2 ;
  RECT 1612.060 0.000 1613.180 1.120 ;
  LAYER metal1 ;
  RECT 1612.060 0.000 1613.180 1.120 ;
 END
END DIA59
PIN DOA59
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1598.420 0.000 1599.540 1.120 ;
  LAYER metal4 ;
  RECT 1598.420 0.000 1599.540 1.120 ;
  LAYER metal3 ;
  RECT 1598.420 0.000 1599.540 1.120 ;
  LAYER metal2 ;
  RECT 1598.420 0.000 1599.540 1.120 ;
  LAYER metal1 ;
  RECT 1598.420 0.000 1599.540 1.120 ;
 END
END DOA59
PIN DIA58
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1585.400 0.000 1586.520 1.120 ;
  LAYER metal4 ;
  RECT 1585.400 0.000 1586.520 1.120 ;
  LAYER metal3 ;
  RECT 1585.400 0.000 1586.520 1.120 ;
  LAYER metal2 ;
  RECT 1585.400 0.000 1586.520 1.120 ;
  LAYER metal1 ;
  RECT 1585.400 0.000 1586.520 1.120 ;
 END
END DIA58
PIN DOA58
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1571.760 0.000 1572.880 1.120 ;
  LAYER metal4 ;
  RECT 1571.760 0.000 1572.880 1.120 ;
  LAYER metal3 ;
  RECT 1571.760 0.000 1572.880 1.120 ;
  LAYER metal2 ;
  RECT 1571.760 0.000 1572.880 1.120 ;
  LAYER metal1 ;
  RECT 1571.760 0.000 1572.880 1.120 ;
 END
END DOA58
PIN DIA57
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1558.120 0.000 1559.240 1.120 ;
  LAYER metal4 ;
  RECT 1558.120 0.000 1559.240 1.120 ;
  LAYER metal3 ;
  RECT 1558.120 0.000 1559.240 1.120 ;
  LAYER metal2 ;
  RECT 1558.120 0.000 1559.240 1.120 ;
  LAYER metal1 ;
  RECT 1558.120 0.000 1559.240 1.120 ;
 END
END DIA57
PIN DOA57
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1545.100 0.000 1546.220 1.120 ;
  LAYER metal4 ;
  RECT 1545.100 0.000 1546.220 1.120 ;
  LAYER metal3 ;
  RECT 1545.100 0.000 1546.220 1.120 ;
  LAYER metal2 ;
  RECT 1545.100 0.000 1546.220 1.120 ;
  LAYER metal1 ;
  RECT 1545.100 0.000 1546.220 1.120 ;
 END
END DOA57
PIN DIA56
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1531.460 0.000 1532.580 1.120 ;
  LAYER metal4 ;
  RECT 1531.460 0.000 1532.580 1.120 ;
  LAYER metal3 ;
  RECT 1531.460 0.000 1532.580 1.120 ;
  LAYER metal2 ;
  RECT 1531.460 0.000 1532.580 1.120 ;
  LAYER metal1 ;
  RECT 1531.460 0.000 1532.580 1.120 ;
 END
END DIA56
PIN DOA56
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1517.820 0.000 1518.940 1.120 ;
  LAYER metal4 ;
  RECT 1517.820 0.000 1518.940 1.120 ;
  LAYER metal3 ;
  RECT 1517.820 0.000 1518.940 1.120 ;
  LAYER metal2 ;
  RECT 1517.820 0.000 1518.940 1.120 ;
  LAYER metal1 ;
  RECT 1517.820 0.000 1518.940 1.120 ;
 END
END DOA56
PIN DIA55
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1504.800 0.000 1505.920 1.120 ;
  LAYER metal4 ;
  RECT 1504.800 0.000 1505.920 1.120 ;
  LAYER metal3 ;
  RECT 1504.800 0.000 1505.920 1.120 ;
  LAYER metal2 ;
  RECT 1504.800 0.000 1505.920 1.120 ;
  LAYER metal1 ;
  RECT 1504.800 0.000 1505.920 1.120 ;
 END
END DIA55
PIN DOA55
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1491.160 0.000 1492.280 1.120 ;
  LAYER metal4 ;
  RECT 1491.160 0.000 1492.280 1.120 ;
  LAYER metal3 ;
  RECT 1491.160 0.000 1492.280 1.120 ;
  LAYER metal2 ;
  RECT 1491.160 0.000 1492.280 1.120 ;
  LAYER metal1 ;
  RECT 1491.160 0.000 1492.280 1.120 ;
 END
END DOA55
PIN DIA54
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1477.520 0.000 1478.640 1.120 ;
  LAYER metal4 ;
  RECT 1477.520 0.000 1478.640 1.120 ;
  LAYER metal3 ;
  RECT 1477.520 0.000 1478.640 1.120 ;
  LAYER metal2 ;
  RECT 1477.520 0.000 1478.640 1.120 ;
  LAYER metal1 ;
  RECT 1477.520 0.000 1478.640 1.120 ;
 END
END DIA54
PIN DOA54
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1464.500 0.000 1465.620 1.120 ;
  LAYER metal4 ;
  RECT 1464.500 0.000 1465.620 1.120 ;
  LAYER metal3 ;
  RECT 1464.500 0.000 1465.620 1.120 ;
  LAYER metal2 ;
  RECT 1464.500 0.000 1465.620 1.120 ;
  LAYER metal1 ;
  RECT 1464.500 0.000 1465.620 1.120 ;
 END
END DOA54
PIN DIA53
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1450.860 0.000 1451.980 1.120 ;
  LAYER metal4 ;
  RECT 1450.860 0.000 1451.980 1.120 ;
  LAYER metal3 ;
  RECT 1450.860 0.000 1451.980 1.120 ;
  LAYER metal2 ;
  RECT 1450.860 0.000 1451.980 1.120 ;
  LAYER metal1 ;
  RECT 1450.860 0.000 1451.980 1.120 ;
 END
END DIA53
PIN DOA53
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1437.220 0.000 1438.340 1.120 ;
  LAYER metal4 ;
  RECT 1437.220 0.000 1438.340 1.120 ;
  LAYER metal3 ;
  RECT 1437.220 0.000 1438.340 1.120 ;
  LAYER metal2 ;
  RECT 1437.220 0.000 1438.340 1.120 ;
  LAYER metal1 ;
  RECT 1437.220 0.000 1438.340 1.120 ;
 END
END DOA53
PIN DIA52
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1424.200 0.000 1425.320 1.120 ;
  LAYER metal4 ;
  RECT 1424.200 0.000 1425.320 1.120 ;
  LAYER metal3 ;
  RECT 1424.200 0.000 1425.320 1.120 ;
  LAYER metal2 ;
  RECT 1424.200 0.000 1425.320 1.120 ;
  LAYER metal1 ;
  RECT 1424.200 0.000 1425.320 1.120 ;
 END
END DIA52
PIN DOA52
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1410.560 0.000 1411.680 1.120 ;
  LAYER metal4 ;
  RECT 1410.560 0.000 1411.680 1.120 ;
  LAYER metal3 ;
  RECT 1410.560 0.000 1411.680 1.120 ;
  LAYER metal2 ;
  RECT 1410.560 0.000 1411.680 1.120 ;
  LAYER metal1 ;
  RECT 1410.560 0.000 1411.680 1.120 ;
 END
END DOA52
PIN DIA51
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1396.920 0.000 1398.040 1.120 ;
  LAYER metal4 ;
  RECT 1396.920 0.000 1398.040 1.120 ;
  LAYER metal3 ;
  RECT 1396.920 0.000 1398.040 1.120 ;
  LAYER metal2 ;
  RECT 1396.920 0.000 1398.040 1.120 ;
  LAYER metal1 ;
  RECT 1396.920 0.000 1398.040 1.120 ;
 END
END DIA51
PIN DOA51
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1383.900 0.000 1385.020 1.120 ;
  LAYER metal4 ;
  RECT 1383.900 0.000 1385.020 1.120 ;
  LAYER metal3 ;
  RECT 1383.900 0.000 1385.020 1.120 ;
  LAYER metal2 ;
  RECT 1383.900 0.000 1385.020 1.120 ;
  LAYER metal1 ;
  RECT 1383.900 0.000 1385.020 1.120 ;
 END
END DOA51
PIN DIA50
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1370.260 0.000 1371.380 1.120 ;
  LAYER metal4 ;
  RECT 1370.260 0.000 1371.380 1.120 ;
  LAYER metal3 ;
  RECT 1370.260 0.000 1371.380 1.120 ;
  LAYER metal2 ;
  RECT 1370.260 0.000 1371.380 1.120 ;
  LAYER metal1 ;
  RECT 1370.260 0.000 1371.380 1.120 ;
 END
END DIA50
PIN DOA50
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1356.620 0.000 1357.740 1.120 ;
  LAYER metal4 ;
  RECT 1356.620 0.000 1357.740 1.120 ;
  LAYER metal3 ;
  RECT 1356.620 0.000 1357.740 1.120 ;
  LAYER metal2 ;
  RECT 1356.620 0.000 1357.740 1.120 ;
  LAYER metal1 ;
  RECT 1356.620 0.000 1357.740 1.120 ;
 END
END DOA50
PIN DIA49
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1343.600 0.000 1344.720 1.120 ;
  LAYER metal4 ;
  RECT 1343.600 0.000 1344.720 1.120 ;
  LAYER metal3 ;
  RECT 1343.600 0.000 1344.720 1.120 ;
  LAYER metal2 ;
  RECT 1343.600 0.000 1344.720 1.120 ;
  LAYER metal1 ;
  RECT 1343.600 0.000 1344.720 1.120 ;
 END
END DIA49
PIN DOA49
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1329.960 0.000 1331.080 1.120 ;
  LAYER metal4 ;
  RECT 1329.960 0.000 1331.080 1.120 ;
  LAYER metal3 ;
  RECT 1329.960 0.000 1331.080 1.120 ;
  LAYER metal2 ;
  RECT 1329.960 0.000 1331.080 1.120 ;
  LAYER metal1 ;
  RECT 1329.960 0.000 1331.080 1.120 ;
 END
END DOA49
PIN DIA48
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1316.320 0.000 1317.440 1.120 ;
  LAYER metal4 ;
  RECT 1316.320 0.000 1317.440 1.120 ;
  LAYER metal3 ;
  RECT 1316.320 0.000 1317.440 1.120 ;
  LAYER metal2 ;
  RECT 1316.320 0.000 1317.440 1.120 ;
  LAYER metal1 ;
  RECT 1316.320 0.000 1317.440 1.120 ;
 END
END DIA48
PIN DOA48
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1302.680 0.000 1303.800 1.120 ;
  LAYER metal4 ;
  RECT 1302.680 0.000 1303.800 1.120 ;
  LAYER metal3 ;
  RECT 1302.680 0.000 1303.800 1.120 ;
  LAYER metal2 ;
  RECT 1302.680 0.000 1303.800 1.120 ;
  LAYER metal1 ;
  RECT 1302.680 0.000 1303.800 1.120 ;
 END
END DOA48
PIN DIA47
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1289.660 0.000 1290.780 1.120 ;
  LAYER metal4 ;
  RECT 1289.660 0.000 1290.780 1.120 ;
  LAYER metal3 ;
  RECT 1289.660 0.000 1290.780 1.120 ;
  LAYER metal2 ;
  RECT 1289.660 0.000 1290.780 1.120 ;
  LAYER metal1 ;
  RECT 1289.660 0.000 1290.780 1.120 ;
 END
END DIA47
PIN DOA47
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1276.020 0.000 1277.140 1.120 ;
  LAYER metal4 ;
  RECT 1276.020 0.000 1277.140 1.120 ;
  LAYER metal3 ;
  RECT 1276.020 0.000 1277.140 1.120 ;
  LAYER metal2 ;
  RECT 1276.020 0.000 1277.140 1.120 ;
  LAYER metal1 ;
  RECT 1276.020 0.000 1277.140 1.120 ;
 END
END DOA47
PIN DIA46
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1262.380 0.000 1263.500 1.120 ;
  LAYER metal4 ;
  RECT 1262.380 0.000 1263.500 1.120 ;
  LAYER metal3 ;
  RECT 1262.380 0.000 1263.500 1.120 ;
  LAYER metal2 ;
  RECT 1262.380 0.000 1263.500 1.120 ;
  LAYER metal1 ;
  RECT 1262.380 0.000 1263.500 1.120 ;
 END
END DIA46
PIN DOA46
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1249.360 0.000 1250.480 1.120 ;
  LAYER metal4 ;
  RECT 1249.360 0.000 1250.480 1.120 ;
  LAYER metal3 ;
  RECT 1249.360 0.000 1250.480 1.120 ;
  LAYER metal2 ;
  RECT 1249.360 0.000 1250.480 1.120 ;
  LAYER metal1 ;
  RECT 1249.360 0.000 1250.480 1.120 ;
 END
END DOA46
PIN DIA45
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1235.720 0.000 1236.840 1.120 ;
  LAYER metal4 ;
  RECT 1235.720 0.000 1236.840 1.120 ;
  LAYER metal3 ;
  RECT 1235.720 0.000 1236.840 1.120 ;
  LAYER metal2 ;
  RECT 1235.720 0.000 1236.840 1.120 ;
  LAYER metal1 ;
  RECT 1235.720 0.000 1236.840 1.120 ;
 END
END DIA45
PIN DOA45
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1222.080 0.000 1223.200 1.120 ;
  LAYER metal4 ;
  RECT 1222.080 0.000 1223.200 1.120 ;
  LAYER metal3 ;
  RECT 1222.080 0.000 1223.200 1.120 ;
  LAYER metal2 ;
  RECT 1222.080 0.000 1223.200 1.120 ;
  LAYER metal1 ;
  RECT 1222.080 0.000 1223.200 1.120 ;
 END
END DOA45
PIN DIA44
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1209.060 0.000 1210.180 1.120 ;
  LAYER metal4 ;
  RECT 1209.060 0.000 1210.180 1.120 ;
  LAYER metal3 ;
  RECT 1209.060 0.000 1210.180 1.120 ;
  LAYER metal2 ;
  RECT 1209.060 0.000 1210.180 1.120 ;
  LAYER metal1 ;
  RECT 1209.060 0.000 1210.180 1.120 ;
 END
END DIA44
PIN DOA44
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1195.420 0.000 1196.540 1.120 ;
  LAYER metal4 ;
  RECT 1195.420 0.000 1196.540 1.120 ;
  LAYER metal3 ;
  RECT 1195.420 0.000 1196.540 1.120 ;
  LAYER metal2 ;
  RECT 1195.420 0.000 1196.540 1.120 ;
  LAYER metal1 ;
  RECT 1195.420 0.000 1196.540 1.120 ;
 END
END DOA44
PIN DIA43
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1181.780 0.000 1182.900 1.120 ;
  LAYER metal4 ;
  RECT 1181.780 0.000 1182.900 1.120 ;
  LAYER metal3 ;
  RECT 1181.780 0.000 1182.900 1.120 ;
  LAYER metal2 ;
  RECT 1181.780 0.000 1182.900 1.120 ;
  LAYER metal1 ;
  RECT 1181.780 0.000 1182.900 1.120 ;
 END
END DIA43
PIN DOA43
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1168.760 0.000 1169.880 1.120 ;
  LAYER metal4 ;
  RECT 1168.760 0.000 1169.880 1.120 ;
  LAYER metal3 ;
  RECT 1168.760 0.000 1169.880 1.120 ;
  LAYER metal2 ;
  RECT 1168.760 0.000 1169.880 1.120 ;
  LAYER metal1 ;
  RECT 1168.760 0.000 1169.880 1.120 ;
 END
END DOA43
PIN DIA42
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1155.120 0.000 1156.240 1.120 ;
  LAYER metal4 ;
  RECT 1155.120 0.000 1156.240 1.120 ;
  LAYER metal3 ;
  RECT 1155.120 0.000 1156.240 1.120 ;
  LAYER metal2 ;
  RECT 1155.120 0.000 1156.240 1.120 ;
  LAYER metal1 ;
  RECT 1155.120 0.000 1156.240 1.120 ;
 END
END DIA42
PIN DOA42
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1141.480 0.000 1142.600 1.120 ;
  LAYER metal4 ;
  RECT 1141.480 0.000 1142.600 1.120 ;
  LAYER metal3 ;
  RECT 1141.480 0.000 1142.600 1.120 ;
  LAYER metal2 ;
  RECT 1141.480 0.000 1142.600 1.120 ;
  LAYER metal1 ;
  RECT 1141.480 0.000 1142.600 1.120 ;
 END
END DOA42
PIN DIA41
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1128.460 0.000 1129.580 1.120 ;
  LAYER metal4 ;
  RECT 1128.460 0.000 1129.580 1.120 ;
  LAYER metal3 ;
  RECT 1128.460 0.000 1129.580 1.120 ;
  LAYER metal2 ;
  RECT 1128.460 0.000 1129.580 1.120 ;
  LAYER metal1 ;
  RECT 1128.460 0.000 1129.580 1.120 ;
 END
END DIA41
PIN DOA41
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1114.820 0.000 1115.940 1.120 ;
  LAYER metal4 ;
  RECT 1114.820 0.000 1115.940 1.120 ;
  LAYER metal3 ;
  RECT 1114.820 0.000 1115.940 1.120 ;
  LAYER metal2 ;
  RECT 1114.820 0.000 1115.940 1.120 ;
  LAYER metal1 ;
  RECT 1114.820 0.000 1115.940 1.120 ;
 END
END DOA41
PIN DIA40
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1101.180 0.000 1102.300 1.120 ;
  LAYER metal4 ;
  RECT 1101.180 0.000 1102.300 1.120 ;
  LAYER metal3 ;
  RECT 1101.180 0.000 1102.300 1.120 ;
  LAYER metal2 ;
  RECT 1101.180 0.000 1102.300 1.120 ;
  LAYER metal1 ;
  RECT 1101.180 0.000 1102.300 1.120 ;
 END
END DIA40
PIN DOA40
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1088.160 0.000 1089.280 1.120 ;
  LAYER metal4 ;
  RECT 1088.160 0.000 1089.280 1.120 ;
  LAYER metal3 ;
  RECT 1088.160 0.000 1089.280 1.120 ;
  LAYER metal2 ;
  RECT 1088.160 0.000 1089.280 1.120 ;
  LAYER metal1 ;
  RECT 1088.160 0.000 1089.280 1.120 ;
 END
END DOA40
PIN DIA39
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1074.520 0.000 1075.640 1.120 ;
  LAYER metal4 ;
  RECT 1074.520 0.000 1075.640 1.120 ;
  LAYER metal3 ;
  RECT 1074.520 0.000 1075.640 1.120 ;
  LAYER metal2 ;
  RECT 1074.520 0.000 1075.640 1.120 ;
  LAYER metal1 ;
  RECT 1074.520 0.000 1075.640 1.120 ;
 END
END DIA39
PIN DOA39
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1060.880 0.000 1062.000 1.120 ;
  LAYER metal4 ;
  RECT 1060.880 0.000 1062.000 1.120 ;
  LAYER metal3 ;
  RECT 1060.880 0.000 1062.000 1.120 ;
  LAYER metal2 ;
  RECT 1060.880 0.000 1062.000 1.120 ;
  LAYER metal1 ;
  RECT 1060.880 0.000 1062.000 1.120 ;
 END
END DOA39
PIN DIA38
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1047.860 0.000 1048.980 1.120 ;
  LAYER metal4 ;
  RECT 1047.860 0.000 1048.980 1.120 ;
  LAYER metal3 ;
  RECT 1047.860 0.000 1048.980 1.120 ;
  LAYER metal2 ;
  RECT 1047.860 0.000 1048.980 1.120 ;
  LAYER metal1 ;
  RECT 1047.860 0.000 1048.980 1.120 ;
 END
END DIA38
PIN DOA38
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1034.220 0.000 1035.340 1.120 ;
  LAYER metal4 ;
  RECT 1034.220 0.000 1035.340 1.120 ;
  LAYER metal3 ;
  RECT 1034.220 0.000 1035.340 1.120 ;
  LAYER metal2 ;
  RECT 1034.220 0.000 1035.340 1.120 ;
  LAYER metal1 ;
  RECT 1034.220 0.000 1035.340 1.120 ;
 END
END DOA38
PIN DIA37
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1020.580 0.000 1021.700 1.120 ;
  LAYER metal4 ;
  RECT 1020.580 0.000 1021.700 1.120 ;
  LAYER metal3 ;
  RECT 1020.580 0.000 1021.700 1.120 ;
  LAYER metal2 ;
  RECT 1020.580 0.000 1021.700 1.120 ;
  LAYER metal1 ;
  RECT 1020.580 0.000 1021.700 1.120 ;
 END
END DIA37
PIN DOA37
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1007.560 0.000 1008.680 1.120 ;
  LAYER metal4 ;
  RECT 1007.560 0.000 1008.680 1.120 ;
  LAYER metal3 ;
  RECT 1007.560 0.000 1008.680 1.120 ;
  LAYER metal2 ;
  RECT 1007.560 0.000 1008.680 1.120 ;
  LAYER metal1 ;
  RECT 1007.560 0.000 1008.680 1.120 ;
 END
END DOA37
PIN DIA36
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 993.920 0.000 995.040 1.120 ;
  LAYER metal4 ;
  RECT 993.920 0.000 995.040 1.120 ;
  LAYER metal3 ;
  RECT 993.920 0.000 995.040 1.120 ;
  LAYER metal2 ;
  RECT 993.920 0.000 995.040 1.120 ;
  LAYER metal1 ;
  RECT 993.920 0.000 995.040 1.120 ;
 END
END DIA36
PIN DOA36
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 980.280 0.000 981.400 1.120 ;
  LAYER metal4 ;
  RECT 980.280 0.000 981.400 1.120 ;
  LAYER metal3 ;
  RECT 980.280 0.000 981.400 1.120 ;
  LAYER metal2 ;
  RECT 980.280 0.000 981.400 1.120 ;
  LAYER metal1 ;
  RECT 980.280 0.000 981.400 1.120 ;
 END
END DOA36
PIN DIA35
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 967.260 0.000 968.380 1.120 ;
  LAYER metal4 ;
  RECT 967.260 0.000 968.380 1.120 ;
  LAYER metal3 ;
  RECT 967.260 0.000 968.380 1.120 ;
  LAYER metal2 ;
  RECT 967.260 0.000 968.380 1.120 ;
  LAYER metal1 ;
  RECT 967.260 0.000 968.380 1.120 ;
 END
END DIA35
PIN DOA35
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 953.620 0.000 954.740 1.120 ;
  LAYER metal4 ;
  RECT 953.620 0.000 954.740 1.120 ;
  LAYER metal3 ;
  RECT 953.620 0.000 954.740 1.120 ;
  LAYER metal2 ;
  RECT 953.620 0.000 954.740 1.120 ;
  LAYER metal1 ;
  RECT 953.620 0.000 954.740 1.120 ;
 END
END DOA35
PIN DIA34
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 939.980 0.000 941.100 1.120 ;
  LAYER metal4 ;
  RECT 939.980 0.000 941.100 1.120 ;
  LAYER metal3 ;
  RECT 939.980 0.000 941.100 1.120 ;
  LAYER metal2 ;
  RECT 939.980 0.000 941.100 1.120 ;
  LAYER metal1 ;
  RECT 939.980 0.000 941.100 1.120 ;
 END
END DIA34
PIN DOA34
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 926.960 0.000 928.080 1.120 ;
  LAYER metal4 ;
  RECT 926.960 0.000 928.080 1.120 ;
  LAYER metal3 ;
  RECT 926.960 0.000 928.080 1.120 ;
  LAYER metal2 ;
  RECT 926.960 0.000 928.080 1.120 ;
  LAYER metal1 ;
  RECT 926.960 0.000 928.080 1.120 ;
 END
END DOA34
PIN DIA33
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 913.320 0.000 914.440 1.120 ;
  LAYER metal4 ;
  RECT 913.320 0.000 914.440 1.120 ;
  LAYER metal3 ;
  RECT 913.320 0.000 914.440 1.120 ;
  LAYER metal2 ;
  RECT 913.320 0.000 914.440 1.120 ;
  LAYER metal1 ;
  RECT 913.320 0.000 914.440 1.120 ;
 END
END DIA33
PIN DOA33
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 899.680 0.000 900.800 1.120 ;
  LAYER metal4 ;
  RECT 899.680 0.000 900.800 1.120 ;
  LAYER metal3 ;
  RECT 899.680 0.000 900.800 1.120 ;
  LAYER metal2 ;
  RECT 899.680 0.000 900.800 1.120 ;
  LAYER metal1 ;
  RECT 899.680 0.000 900.800 1.120 ;
 END
END DOA33
PIN DIA32
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 886.040 0.000 887.160 1.120 ;
  LAYER metal4 ;
  RECT 886.040 0.000 887.160 1.120 ;
  LAYER metal3 ;
  RECT 886.040 0.000 887.160 1.120 ;
  LAYER metal2 ;
  RECT 886.040 0.000 887.160 1.120 ;
  LAYER metal1 ;
  RECT 886.040 0.000 887.160 1.120 ;
 END
END DIA32
PIN DOA32
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 873.020 0.000 874.140 1.120 ;
  LAYER metal4 ;
  RECT 873.020 0.000 874.140 1.120 ;
  LAYER metal3 ;
  RECT 873.020 0.000 874.140 1.120 ;
  LAYER metal2 ;
  RECT 873.020 0.000 874.140 1.120 ;
  LAYER metal1 ;
  RECT 873.020 0.000 874.140 1.120 ;
 END
END DOA32
PIN DIA31
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 859.380 0.000 860.500 1.120 ;
  LAYER metal4 ;
  RECT 859.380 0.000 860.500 1.120 ;
  LAYER metal3 ;
  RECT 859.380 0.000 860.500 1.120 ;
  LAYER metal2 ;
  RECT 859.380 0.000 860.500 1.120 ;
  LAYER metal1 ;
  RECT 859.380 0.000 860.500 1.120 ;
 END
END DIA31
PIN DOA31
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 845.740 0.000 846.860 1.120 ;
  LAYER metal4 ;
  RECT 845.740 0.000 846.860 1.120 ;
  LAYER metal3 ;
  RECT 845.740 0.000 846.860 1.120 ;
  LAYER metal2 ;
  RECT 845.740 0.000 846.860 1.120 ;
  LAYER metal1 ;
  RECT 845.740 0.000 846.860 1.120 ;
 END
END DOA31
PIN DIA30
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 832.720 0.000 833.840 1.120 ;
  LAYER metal4 ;
  RECT 832.720 0.000 833.840 1.120 ;
  LAYER metal3 ;
  RECT 832.720 0.000 833.840 1.120 ;
  LAYER metal2 ;
  RECT 832.720 0.000 833.840 1.120 ;
  LAYER metal1 ;
  RECT 832.720 0.000 833.840 1.120 ;
 END
END DIA30
PIN DOA30
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 819.080 0.000 820.200 1.120 ;
  LAYER metal4 ;
  RECT 819.080 0.000 820.200 1.120 ;
  LAYER metal3 ;
  RECT 819.080 0.000 820.200 1.120 ;
  LAYER metal2 ;
  RECT 819.080 0.000 820.200 1.120 ;
  LAYER metal1 ;
  RECT 819.080 0.000 820.200 1.120 ;
 END
END DOA30
PIN DIA29
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 805.440 0.000 806.560 1.120 ;
  LAYER metal4 ;
  RECT 805.440 0.000 806.560 1.120 ;
  LAYER metal3 ;
  RECT 805.440 0.000 806.560 1.120 ;
  LAYER metal2 ;
  RECT 805.440 0.000 806.560 1.120 ;
  LAYER metal1 ;
  RECT 805.440 0.000 806.560 1.120 ;
 END
END DIA29
PIN DOA29
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 792.420 0.000 793.540 1.120 ;
  LAYER metal4 ;
  RECT 792.420 0.000 793.540 1.120 ;
  LAYER metal3 ;
  RECT 792.420 0.000 793.540 1.120 ;
  LAYER metal2 ;
  RECT 792.420 0.000 793.540 1.120 ;
  LAYER metal1 ;
  RECT 792.420 0.000 793.540 1.120 ;
 END
END DOA29
PIN DIA28
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 778.780 0.000 779.900 1.120 ;
  LAYER metal4 ;
  RECT 778.780 0.000 779.900 1.120 ;
  LAYER metal3 ;
  RECT 778.780 0.000 779.900 1.120 ;
  LAYER metal2 ;
  RECT 778.780 0.000 779.900 1.120 ;
  LAYER metal1 ;
  RECT 778.780 0.000 779.900 1.120 ;
 END
END DIA28
PIN DOA28
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 765.140 0.000 766.260 1.120 ;
  LAYER metal4 ;
  RECT 765.140 0.000 766.260 1.120 ;
  LAYER metal3 ;
  RECT 765.140 0.000 766.260 1.120 ;
  LAYER metal2 ;
  RECT 765.140 0.000 766.260 1.120 ;
  LAYER metal1 ;
  RECT 765.140 0.000 766.260 1.120 ;
 END
END DOA28
PIN DIA27
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 752.120 0.000 753.240 1.120 ;
  LAYER metal4 ;
  RECT 752.120 0.000 753.240 1.120 ;
  LAYER metal3 ;
  RECT 752.120 0.000 753.240 1.120 ;
  LAYER metal2 ;
  RECT 752.120 0.000 753.240 1.120 ;
  LAYER metal1 ;
  RECT 752.120 0.000 753.240 1.120 ;
 END
END DIA27
PIN DOA27
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 738.480 0.000 739.600 1.120 ;
  LAYER metal4 ;
  RECT 738.480 0.000 739.600 1.120 ;
  LAYER metal3 ;
  RECT 738.480 0.000 739.600 1.120 ;
  LAYER metal2 ;
  RECT 738.480 0.000 739.600 1.120 ;
  LAYER metal1 ;
  RECT 738.480 0.000 739.600 1.120 ;
 END
END DOA27
PIN DIA26
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 724.840 0.000 725.960 1.120 ;
  LAYER metal4 ;
  RECT 724.840 0.000 725.960 1.120 ;
  LAYER metal3 ;
  RECT 724.840 0.000 725.960 1.120 ;
  LAYER metal2 ;
  RECT 724.840 0.000 725.960 1.120 ;
  LAYER metal1 ;
  RECT 724.840 0.000 725.960 1.120 ;
 END
END DIA26
PIN DOA26
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 711.820 0.000 712.940 1.120 ;
  LAYER metal4 ;
  RECT 711.820 0.000 712.940 1.120 ;
  LAYER metal3 ;
  RECT 711.820 0.000 712.940 1.120 ;
  LAYER metal2 ;
  RECT 711.820 0.000 712.940 1.120 ;
  LAYER metal1 ;
  RECT 711.820 0.000 712.940 1.120 ;
 END
END DOA26
PIN DIA25
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 698.180 0.000 699.300 1.120 ;
  LAYER metal4 ;
  RECT 698.180 0.000 699.300 1.120 ;
  LAYER metal3 ;
  RECT 698.180 0.000 699.300 1.120 ;
  LAYER metal2 ;
  RECT 698.180 0.000 699.300 1.120 ;
  LAYER metal1 ;
  RECT 698.180 0.000 699.300 1.120 ;
 END
END DIA25
PIN DOA25
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 684.540 0.000 685.660 1.120 ;
  LAYER metal4 ;
  RECT 684.540 0.000 685.660 1.120 ;
  LAYER metal3 ;
  RECT 684.540 0.000 685.660 1.120 ;
  LAYER metal2 ;
  RECT 684.540 0.000 685.660 1.120 ;
  LAYER metal1 ;
  RECT 684.540 0.000 685.660 1.120 ;
 END
END DOA25
PIN DIA24
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 671.520 0.000 672.640 1.120 ;
  LAYER metal4 ;
  RECT 671.520 0.000 672.640 1.120 ;
  LAYER metal3 ;
  RECT 671.520 0.000 672.640 1.120 ;
  LAYER metal2 ;
  RECT 671.520 0.000 672.640 1.120 ;
  LAYER metal1 ;
  RECT 671.520 0.000 672.640 1.120 ;
 END
END DIA24
PIN DOA24
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 657.880 0.000 659.000 1.120 ;
  LAYER metal4 ;
  RECT 657.880 0.000 659.000 1.120 ;
  LAYER metal3 ;
  RECT 657.880 0.000 659.000 1.120 ;
  LAYER metal2 ;
  RECT 657.880 0.000 659.000 1.120 ;
  LAYER metal1 ;
  RECT 657.880 0.000 659.000 1.120 ;
 END
END DOA24
PIN DIA23
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 644.240 0.000 645.360 1.120 ;
  LAYER metal4 ;
  RECT 644.240 0.000 645.360 1.120 ;
  LAYER metal3 ;
  RECT 644.240 0.000 645.360 1.120 ;
  LAYER metal2 ;
  RECT 644.240 0.000 645.360 1.120 ;
  LAYER metal1 ;
  RECT 644.240 0.000 645.360 1.120 ;
 END
END DIA23
PIN DOA23
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 631.220 0.000 632.340 1.120 ;
  LAYER metal4 ;
  RECT 631.220 0.000 632.340 1.120 ;
  LAYER metal3 ;
  RECT 631.220 0.000 632.340 1.120 ;
  LAYER metal2 ;
  RECT 631.220 0.000 632.340 1.120 ;
  LAYER metal1 ;
  RECT 631.220 0.000 632.340 1.120 ;
 END
END DOA23
PIN DIA22
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 617.580 0.000 618.700 1.120 ;
  LAYER metal4 ;
  RECT 617.580 0.000 618.700 1.120 ;
  LAYER metal3 ;
  RECT 617.580 0.000 618.700 1.120 ;
  LAYER metal2 ;
  RECT 617.580 0.000 618.700 1.120 ;
  LAYER metal1 ;
  RECT 617.580 0.000 618.700 1.120 ;
 END
END DIA22
PIN DOA22
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 603.940 0.000 605.060 1.120 ;
  LAYER metal4 ;
  RECT 603.940 0.000 605.060 1.120 ;
  LAYER metal3 ;
  RECT 603.940 0.000 605.060 1.120 ;
  LAYER metal2 ;
  RECT 603.940 0.000 605.060 1.120 ;
  LAYER metal1 ;
  RECT 603.940 0.000 605.060 1.120 ;
 END
END DOA22
PIN DIA21
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 590.920 0.000 592.040 1.120 ;
  LAYER metal4 ;
  RECT 590.920 0.000 592.040 1.120 ;
  LAYER metal3 ;
  RECT 590.920 0.000 592.040 1.120 ;
  LAYER metal2 ;
  RECT 590.920 0.000 592.040 1.120 ;
  LAYER metal1 ;
  RECT 590.920 0.000 592.040 1.120 ;
 END
END DIA21
PIN DOA21
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 577.280 0.000 578.400 1.120 ;
  LAYER metal4 ;
  RECT 577.280 0.000 578.400 1.120 ;
  LAYER metal3 ;
  RECT 577.280 0.000 578.400 1.120 ;
  LAYER metal2 ;
  RECT 577.280 0.000 578.400 1.120 ;
  LAYER metal1 ;
  RECT 577.280 0.000 578.400 1.120 ;
 END
END DOA21
PIN DIA20
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 563.640 0.000 564.760 1.120 ;
  LAYER metal4 ;
  RECT 563.640 0.000 564.760 1.120 ;
  LAYER metal3 ;
  RECT 563.640 0.000 564.760 1.120 ;
  LAYER metal2 ;
  RECT 563.640 0.000 564.760 1.120 ;
  LAYER metal1 ;
  RECT 563.640 0.000 564.760 1.120 ;
 END
END DIA20
PIN DOA20
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 550.620 0.000 551.740 1.120 ;
  LAYER metal4 ;
  RECT 550.620 0.000 551.740 1.120 ;
  LAYER metal3 ;
  RECT 550.620 0.000 551.740 1.120 ;
  LAYER metal2 ;
  RECT 550.620 0.000 551.740 1.120 ;
  LAYER metal1 ;
  RECT 550.620 0.000 551.740 1.120 ;
 END
END DOA20
PIN DIA19
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 536.980 0.000 538.100 1.120 ;
  LAYER metal4 ;
  RECT 536.980 0.000 538.100 1.120 ;
  LAYER metal3 ;
  RECT 536.980 0.000 538.100 1.120 ;
  LAYER metal2 ;
  RECT 536.980 0.000 538.100 1.120 ;
  LAYER metal1 ;
  RECT 536.980 0.000 538.100 1.120 ;
 END
END DIA19
PIN DOA19
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 523.340 0.000 524.460 1.120 ;
  LAYER metal4 ;
  RECT 523.340 0.000 524.460 1.120 ;
  LAYER metal3 ;
  RECT 523.340 0.000 524.460 1.120 ;
  LAYER metal2 ;
  RECT 523.340 0.000 524.460 1.120 ;
  LAYER metal1 ;
  RECT 523.340 0.000 524.460 1.120 ;
 END
END DOA19
PIN DIA18
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 510.320 0.000 511.440 1.120 ;
  LAYER metal4 ;
  RECT 510.320 0.000 511.440 1.120 ;
  LAYER metal3 ;
  RECT 510.320 0.000 511.440 1.120 ;
  LAYER metal2 ;
  RECT 510.320 0.000 511.440 1.120 ;
  LAYER metal1 ;
  RECT 510.320 0.000 511.440 1.120 ;
 END
END DIA18
PIN DOA18
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 496.680 0.000 497.800 1.120 ;
  LAYER metal4 ;
  RECT 496.680 0.000 497.800 1.120 ;
  LAYER metal3 ;
  RECT 496.680 0.000 497.800 1.120 ;
  LAYER metal2 ;
  RECT 496.680 0.000 497.800 1.120 ;
  LAYER metal1 ;
  RECT 496.680 0.000 497.800 1.120 ;
 END
END DOA18
PIN DIA17
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 483.040 0.000 484.160 1.120 ;
  LAYER metal4 ;
  RECT 483.040 0.000 484.160 1.120 ;
  LAYER metal3 ;
  RECT 483.040 0.000 484.160 1.120 ;
  LAYER metal2 ;
  RECT 483.040 0.000 484.160 1.120 ;
  LAYER metal1 ;
  RECT 483.040 0.000 484.160 1.120 ;
 END
END DIA17
PIN DOA17
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 469.400 0.000 470.520 1.120 ;
  LAYER metal4 ;
  RECT 469.400 0.000 470.520 1.120 ;
  LAYER metal3 ;
  RECT 469.400 0.000 470.520 1.120 ;
  LAYER metal2 ;
  RECT 469.400 0.000 470.520 1.120 ;
  LAYER metal1 ;
  RECT 469.400 0.000 470.520 1.120 ;
 END
END DOA17
PIN DIA16
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 456.380 0.000 457.500 1.120 ;
  LAYER metal4 ;
  RECT 456.380 0.000 457.500 1.120 ;
  LAYER metal3 ;
  RECT 456.380 0.000 457.500 1.120 ;
  LAYER metal2 ;
  RECT 456.380 0.000 457.500 1.120 ;
  LAYER metal1 ;
  RECT 456.380 0.000 457.500 1.120 ;
 END
END DIA16
PIN DOA16
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 442.740 0.000 443.860 1.120 ;
  LAYER metal4 ;
  RECT 442.740 0.000 443.860 1.120 ;
  LAYER metal3 ;
  RECT 442.740 0.000 443.860 1.120 ;
  LAYER metal2 ;
  RECT 442.740 0.000 443.860 1.120 ;
  LAYER metal1 ;
  RECT 442.740 0.000 443.860 1.120 ;
 END
END DOA16
PIN DIA15
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER metal4 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER metal3 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER metal2 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER metal1 ;
  RECT 429.100 0.000 430.220 1.120 ;
 END
END DIA15
PIN DOA15
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 416.080 0.000 417.200 1.120 ;
  LAYER metal4 ;
  RECT 416.080 0.000 417.200 1.120 ;
  LAYER metal3 ;
  RECT 416.080 0.000 417.200 1.120 ;
  LAYER metal2 ;
  RECT 416.080 0.000 417.200 1.120 ;
  LAYER metal1 ;
  RECT 416.080 0.000 417.200 1.120 ;
 END
END DOA15
PIN DIA14
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER metal4 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER metal3 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER metal2 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER metal1 ;
  RECT 402.440 0.000 403.560 1.120 ;
 END
END DIA14
PIN DOA14
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 388.800 0.000 389.920 1.120 ;
  LAYER metal4 ;
  RECT 388.800 0.000 389.920 1.120 ;
  LAYER metal3 ;
  RECT 388.800 0.000 389.920 1.120 ;
  LAYER metal2 ;
  RECT 388.800 0.000 389.920 1.120 ;
  LAYER metal1 ;
  RECT 388.800 0.000 389.920 1.120 ;
 END
END DOA14
PIN DIA13
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 375.780 0.000 376.900 1.120 ;
  LAYER metal4 ;
  RECT 375.780 0.000 376.900 1.120 ;
  LAYER metal3 ;
  RECT 375.780 0.000 376.900 1.120 ;
  LAYER metal2 ;
  RECT 375.780 0.000 376.900 1.120 ;
  LAYER metal1 ;
  RECT 375.780 0.000 376.900 1.120 ;
 END
END DIA13
PIN DOA13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 362.140 0.000 363.260 1.120 ;
  LAYER metal4 ;
  RECT 362.140 0.000 363.260 1.120 ;
  LAYER metal3 ;
  RECT 362.140 0.000 363.260 1.120 ;
  LAYER metal2 ;
  RECT 362.140 0.000 363.260 1.120 ;
  LAYER metal1 ;
  RECT 362.140 0.000 363.260 1.120 ;
 END
END DOA13
PIN DIA12
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 348.500 0.000 349.620 1.120 ;
  LAYER metal4 ;
  RECT 348.500 0.000 349.620 1.120 ;
  LAYER metal3 ;
  RECT 348.500 0.000 349.620 1.120 ;
  LAYER metal2 ;
  RECT 348.500 0.000 349.620 1.120 ;
  LAYER metal1 ;
  RECT 348.500 0.000 349.620 1.120 ;
 END
END DIA12
PIN DOA12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 335.480 0.000 336.600 1.120 ;
  LAYER metal4 ;
  RECT 335.480 0.000 336.600 1.120 ;
  LAYER metal3 ;
  RECT 335.480 0.000 336.600 1.120 ;
  LAYER metal2 ;
  RECT 335.480 0.000 336.600 1.120 ;
  LAYER metal1 ;
  RECT 335.480 0.000 336.600 1.120 ;
 END
END DOA12
PIN DIA11
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 321.840 0.000 322.960 1.120 ;
  LAYER metal4 ;
  RECT 321.840 0.000 322.960 1.120 ;
  LAYER metal3 ;
  RECT 321.840 0.000 322.960 1.120 ;
  LAYER metal2 ;
  RECT 321.840 0.000 322.960 1.120 ;
  LAYER metal1 ;
  RECT 321.840 0.000 322.960 1.120 ;
 END
END DIA11
PIN DOA11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 308.200 0.000 309.320 1.120 ;
  LAYER metal4 ;
  RECT 308.200 0.000 309.320 1.120 ;
  LAYER metal3 ;
  RECT 308.200 0.000 309.320 1.120 ;
  LAYER metal2 ;
  RECT 308.200 0.000 309.320 1.120 ;
  LAYER metal1 ;
  RECT 308.200 0.000 309.320 1.120 ;
 END
END DOA11
PIN DIA10
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 295.180 0.000 296.300 1.120 ;
  LAYER metal4 ;
  RECT 295.180 0.000 296.300 1.120 ;
  LAYER metal3 ;
  RECT 295.180 0.000 296.300 1.120 ;
  LAYER metal2 ;
  RECT 295.180 0.000 296.300 1.120 ;
  LAYER metal1 ;
  RECT 295.180 0.000 296.300 1.120 ;
 END
END DIA10
PIN DOA10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 281.540 0.000 282.660 1.120 ;
  LAYER metal4 ;
  RECT 281.540 0.000 282.660 1.120 ;
  LAYER metal3 ;
  RECT 281.540 0.000 282.660 1.120 ;
  LAYER metal2 ;
  RECT 281.540 0.000 282.660 1.120 ;
  LAYER metal1 ;
  RECT 281.540 0.000 282.660 1.120 ;
 END
END DOA10
PIN DIA9
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER metal4 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER metal3 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER metal2 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER metal1 ;
  RECT 267.900 0.000 269.020 1.120 ;
 END
END DIA9
PIN DOA9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER metal4 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER metal3 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER metal2 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER metal1 ;
  RECT 254.880 0.000 256.000 1.120 ;
 END
END DOA9
PIN DIA8
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER metal4 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER metal3 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER metal2 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER metal1 ;
  RECT 241.240 0.000 242.360 1.120 ;
 END
END DIA8
PIN DOA8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 227.600 0.000 228.720 1.120 ;
  LAYER metal4 ;
  RECT 227.600 0.000 228.720 1.120 ;
  LAYER metal3 ;
  RECT 227.600 0.000 228.720 1.120 ;
  LAYER metal2 ;
  RECT 227.600 0.000 228.720 1.120 ;
  LAYER metal1 ;
  RECT 227.600 0.000 228.720 1.120 ;
 END
END DOA8
PIN DIA7
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 214.580 0.000 215.700 1.120 ;
  LAYER metal4 ;
  RECT 214.580 0.000 215.700 1.120 ;
  LAYER metal3 ;
  RECT 214.580 0.000 215.700 1.120 ;
  LAYER metal2 ;
  RECT 214.580 0.000 215.700 1.120 ;
  LAYER metal1 ;
  RECT 214.580 0.000 215.700 1.120 ;
 END
END DIA7
PIN DOA7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 200.940 0.000 202.060 1.120 ;
  LAYER metal4 ;
  RECT 200.940 0.000 202.060 1.120 ;
  LAYER metal3 ;
  RECT 200.940 0.000 202.060 1.120 ;
  LAYER metal2 ;
  RECT 200.940 0.000 202.060 1.120 ;
  LAYER metal1 ;
  RECT 200.940 0.000 202.060 1.120 ;
 END
END DOA7
PIN DIA6
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER metal4 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER metal3 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER metal2 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER metal1 ;
  RECT 187.300 0.000 188.420 1.120 ;
 END
END DIA6
PIN DOA6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 174.280 0.000 175.400 1.120 ;
  LAYER metal4 ;
  RECT 174.280 0.000 175.400 1.120 ;
  LAYER metal3 ;
  RECT 174.280 0.000 175.400 1.120 ;
  LAYER metal2 ;
  RECT 174.280 0.000 175.400 1.120 ;
  LAYER metal1 ;
  RECT 174.280 0.000 175.400 1.120 ;
 END
END DOA6
PIN DIA5
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 160.640 0.000 161.760 1.120 ;
  LAYER metal4 ;
  RECT 160.640 0.000 161.760 1.120 ;
  LAYER metal3 ;
  RECT 160.640 0.000 161.760 1.120 ;
  LAYER metal2 ;
  RECT 160.640 0.000 161.760 1.120 ;
  LAYER metal1 ;
  RECT 160.640 0.000 161.760 1.120 ;
 END
END DIA5
PIN DOA5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 147.000 0.000 148.120 1.120 ;
  LAYER metal4 ;
  RECT 147.000 0.000 148.120 1.120 ;
  LAYER metal3 ;
  RECT 147.000 0.000 148.120 1.120 ;
  LAYER metal2 ;
  RECT 147.000 0.000 148.120 1.120 ;
  LAYER metal1 ;
  RECT 147.000 0.000 148.120 1.120 ;
 END
END DOA5
PIN DIA4
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 133.980 0.000 135.100 1.120 ;
  LAYER metal4 ;
  RECT 133.980 0.000 135.100 1.120 ;
  LAYER metal3 ;
  RECT 133.980 0.000 135.100 1.120 ;
  LAYER metal2 ;
  RECT 133.980 0.000 135.100 1.120 ;
  LAYER metal1 ;
  RECT 133.980 0.000 135.100 1.120 ;
 END
END DIA4
PIN DOA4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 120.340 0.000 121.460 1.120 ;
  LAYER metal4 ;
  RECT 120.340 0.000 121.460 1.120 ;
  LAYER metal3 ;
  RECT 120.340 0.000 121.460 1.120 ;
  LAYER metal2 ;
  RECT 120.340 0.000 121.460 1.120 ;
  LAYER metal1 ;
  RECT 120.340 0.000 121.460 1.120 ;
 END
END DOA4
PIN DIA3
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal4 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal3 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal2 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal1 ;
  RECT 106.700 0.000 107.820 1.120 ;
 END
END DIA3
PIN DOA3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 93.680 0.000 94.800 1.120 ;
  LAYER metal4 ;
  RECT 93.680 0.000 94.800 1.120 ;
  LAYER metal3 ;
  RECT 93.680 0.000 94.800 1.120 ;
  LAYER metal2 ;
  RECT 93.680 0.000 94.800 1.120 ;
  LAYER metal1 ;
  RECT 93.680 0.000 94.800 1.120 ;
 END
END DOA3
PIN DIA2
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 80.040 0.000 81.160 1.120 ;
  LAYER metal4 ;
  RECT 80.040 0.000 81.160 1.120 ;
  LAYER metal3 ;
  RECT 80.040 0.000 81.160 1.120 ;
  LAYER metal2 ;
  RECT 80.040 0.000 81.160 1.120 ;
  LAYER metal1 ;
  RECT 80.040 0.000 81.160 1.120 ;
 END
END DIA2
PIN DOA2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 66.400 0.000 67.520 1.120 ;
  LAYER metal4 ;
  RECT 66.400 0.000 67.520 1.120 ;
  LAYER metal3 ;
  RECT 66.400 0.000 67.520 1.120 ;
  LAYER metal2 ;
  RECT 66.400 0.000 67.520 1.120 ;
  LAYER metal1 ;
  RECT 66.400 0.000 67.520 1.120 ;
 END
END DOA2
PIN DIA1
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 52.760 0.000 53.880 1.120 ;
  LAYER metal4 ;
  RECT 52.760 0.000 53.880 1.120 ;
  LAYER metal3 ;
  RECT 52.760 0.000 53.880 1.120 ;
  LAYER metal2 ;
  RECT 52.760 0.000 53.880 1.120 ;
  LAYER metal1 ;
  RECT 52.760 0.000 53.880 1.120 ;
 END
END DIA1
PIN DOA1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 39.740 0.000 40.860 1.120 ;
  LAYER metal4 ;
  RECT 39.740 0.000 40.860 1.120 ;
  LAYER metal3 ;
  RECT 39.740 0.000 40.860 1.120 ;
  LAYER metal2 ;
  RECT 39.740 0.000 40.860 1.120 ;
  LAYER metal1 ;
  RECT 39.740 0.000 40.860 1.120 ;
 END
END DOA1
PIN DIA0
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 26.100 0.000 27.220 1.120 ;
  LAYER metal4 ;
  RECT 26.100 0.000 27.220 1.120 ;
  LAYER metal3 ;
  RECT 26.100 0.000 27.220 1.120 ;
  LAYER metal2 ;
  RECT 26.100 0.000 27.220 1.120 ;
  LAYER metal1 ;
  RECT 26.100 0.000 27.220 1.120 ;
 END
END DIA0
PIN DOA0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 12.460 0.000 13.580 1.120 ;
  LAYER metal4 ;
  RECT 12.460 0.000 13.580 1.120 ;
  LAYER metal3 ;
  RECT 12.460 0.000 13.580 1.120 ;
  LAYER metal2 ;
  RECT 12.460 0.000 13.580 1.120 ;
  LAYER metal1 ;
  RECT 12.460 0.000 13.580 1.120 ;
 END
END DOA0
OBS
  LAYER metal1 SPACING 0.280 ;
  RECT 0.000 0.140 3596.000 501.620 ;
  LAYER metal2 SPACING 0.320 ;
  RECT 0.000 0.140 3596.000 501.620 ;
  LAYER metal3 SPACING 0.320 ;
  RECT 0.000 0.140 3596.000 501.620 ;
  LAYER metal4 SPACING 0.600 ;
  RECT 0.000 0.140 3596.000 501.620 ;
  LAYER via ;
  RECT 0.000 0.140 3596.000 501.620 ;
  LAYER via2 ;
  RECT 0.000 0.140 3596.000 501.620 ;
  LAYER via3 ;
  RECT 0.000 0.140 3596.000 501.620 ;
END
END layer1_sram
END LIBRARY



