# 
#              Synchronous Dual Port SRAM Compiler 
# 
#                    UMC 0.18um Generic Logic Process 
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2009 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http://www.faraday-tech.com/
#   
#       Module Name      : layer4_sram
#       Words            : 144
#       Bits             : 128
#       Byte-Write       : 1
#       Aspect Ratio     : 1
#       Output Loading   : 0.5  (pf)
#       Data Slew        : 2.0  (ns)
#       CK Slew          : 2.0  (ns)
#       Power Ring Width : 2  (um)
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSA0M_A
#       Memaker          : 200901.2.1
#       Date             : 2021/01/15 13:26:42
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO layer4_sram
CLASS BLOCK ;
FOREIGN layer4_sram 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 3571.820 BY 210.000 ;
SYMMETRY x y r90 ;
SITE core ;
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal5 ;
  RECT 3570.700 199.700 3571.820 202.940 ;
  LAYER metal4 ;
  RECT 3570.700 199.700 3571.820 202.940 ;
  LAYER metal3 ;
  RECT 3570.700 199.700 3571.820 202.940 ;
  LAYER metal2 ;
  RECT 3570.700 199.700 3571.820 202.940 ;
  LAYER metal1 ;
  RECT 3570.700 199.700 3571.820 202.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.700 191.860 3571.820 195.100 ;
  LAYER metal4 ;
  RECT 3570.700 191.860 3571.820 195.100 ;
  LAYER metal3 ;
  RECT 3570.700 191.860 3571.820 195.100 ;
  LAYER metal2 ;
  RECT 3570.700 191.860 3571.820 195.100 ;
  LAYER metal1 ;
  RECT 3570.700 191.860 3571.820 195.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.700 184.020 3571.820 187.260 ;
  LAYER metal4 ;
  RECT 3570.700 184.020 3571.820 187.260 ;
  LAYER metal3 ;
  RECT 3570.700 184.020 3571.820 187.260 ;
  LAYER metal2 ;
  RECT 3570.700 184.020 3571.820 187.260 ;
  LAYER metal1 ;
  RECT 3570.700 184.020 3571.820 187.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.700 176.180 3571.820 179.420 ;
  LAYER metal4 ;
  RECT 3570.700 176.180 3571.820 179.420 ;
  LAYER metal3 ;
  RECT 3570.700 176.180 3571.820 179.420 ;
  LAYER metal2 ;
  RECT 3570.700 176.180 3571.820 179.420 ;
  LAYER metal1 ;
  RECT 3570.700 176.180 3571.820 179.420 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.700 168.340 3571.820 171.580 ;
  LAYER metal4 ;
  RECT 3570.700 168.340 3571.820 171.580 ;
  LAYER metal3 ;
  RECT 3570.700 168.340 3571.820 171.580 ;
  LAYER metal2 ;
  RECT 3570.700 168.340 3571.820 171.580 ;
  LAYER metal1 ;
  RECT 3570.700 168.340 3571.820 171.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.700 129.140 3571.820 132.380 ;
  LAYER metal4 ;
  RECT 3570.700 129.140 3571.820 132.380 ;
  LAYER metal3 ;
  RECT 3570.700 129.140 3571.820 132.380 ;
  LAYER metal2 ;
  RECT 3570.700 129.140 3571.820 132.380 ;
  LAYER metal1 ;
  RECT 3570.700 129.140 3571.820 132.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.700 121.300 3571.820 124.540 ;
  LAYER metal4 ;
  RECT 3570.700 121.300 3571.820 124.540 ;
  LAYER metal3 ;
  RECT 3570.700 121.300 3571.820 124.540 ;
  LAYER metal2 ;
  RECT 3570.700 121.300 3571.820 124.540 ;
  LAYER metal1 ;
  RECT 3570.700 121.300 3571.820 124.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.700 113.460 3571.820 116.700 ;
  LAYER metal4 ;
  RECT 3570.700 113.460 3571.820 116.700 ;
  LAYER metal3 ;
  RECT 3570.700 113.460 3571.820 116.700 ;
  LAYER metal2 ;
  RECT 3570.700 113.460 3571.820 116.700 ;
  LAYER metal1 ;
  RECT 3570.700 113.460 3571.820 116.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.700 105.620 3571.820 108.860 ;
  LAYER metal4 ;
  RECT 3570.700 105.620 3571.820 108.860 ;
  LAYER metal3 ;
  RECT 3570.700 105.620 3571.820 108.860 ;
  LAYER metal2 ;
  RECT 3570.700 105.620 3571.820 108.860 ;
  LAYER metal1 ;
  RECT 3570.700 105.620 3571.820 108.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.700 97.780 3571.820 101.020 ;
  LAYER metal4 ;
  RECT 3570.700 97.780 3571.820 101.020 ;
  LAYER metal3 ;
  RECT 3570.700 97.780 3571.820 101.020 ;
  LAYER metal2 ;
  RECT 3570.700 97.780 3571.820 101.020 ;
  LAYER metal1 ;
  RECT 3570.700 97.780 3571.820 101.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.700 89.940 3571.820 93.180 ;
  LAYER metal4 ;
  RECT 3570.700 89.940 3571.820 93.180 ;
  LAYER metal3 ;
  RECT 3570.700 89.940 3571.820 93.180 ;
  LAYER metal2 ;
  RECT 3570.700 89.940 3571.820 93.180 ;
  LAYER metal1 ;
  RECT 3570.700 89.940 3571.820 93.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.700 50.740 3571.820 53.980 ;
  LAYER metal4 ;
  RECT 3570.700 50.740 3571.820 53.980 ;
  LAYER metal3 ;
  RECT 3570.700 50.740 3571.820 53.980 ;
  LAYER metal2 ;
  RECT 3570.700 50.740 3571.820 53.980 ;
  LAYER metal1 ;
  RECT 3570.700 50.740 3571.820 53.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.700 42.900 3571.820 46.140 ;
  LAYER metal4 ;
  RECT 3570.700 42.900 3571.820 46.140 ;
  LAYER metal3 ;
  RECT 3570.700 42.900 3571.820 46.140 ;
  LAYER metal2 ;
  RECT 3570.700 42.900 3571.820 46.140 ;
  LAYER metal1 ;
  RECT 3570.700 42.900 3571.820 46.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.700 35.060 3571.820 38.300 ;
  LAYER metal4 ;
  RECT 3570.700 35.060 3571.820 38.300 ;
  LAYER metal3 ;
  RECT 3570.700 35.060 3571.820 38.300 ;
  LAYER metal2 ;
  RECT 3570.700 35.060 3571.820 38.300 ;
  LAYER metal1 ;
  RECT 3570.700 35.060 3571.820 38.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.700 27.220 3571.820 30.460 ;
  LAYER metal4 ;
  RECT 3570.700 27.220 3571.820 30.460 ;
  LAYER metal3 ;
  RECT 3570.700 27.220 3571.820 30.460 ;
  LAYER metal2 ;
  RECT 3570.700 27.220 3571.820 30.460 ;
  LAYER metal1 ;
  RECT 3570.700 27.220 3571.820 30.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.700 19.380 3571.820 22.620 ;
  LAYER metal4 ;
  RECT 3570.700 19.380 3571.820 22.620 ;
  LAYER metal3 ;
  RECT 3570.700 19.380 3571.820 22.620 ;
  LAYER metal2 ;
  RECT 3570.700 19.380 3571.820 22.620 ;
  LAYER metal1 ;
  RECT 3570.700 19.380 3571.820 22.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.700 11.540 3571.820 14.780 ;
  LAYER metal4 ;
  RECT 3570.700 11.540 3571.820 14.780 ;
  LAYER metal3 ;
  RECT 3570.700 11.540 3571.820 14.780 ;
  LAYER metal2 ;
  RECT 3570.700 11.540 3571.820 14.780 ;
  LAYER metal1 ;
  RECT 3570.700 11.540 3571.820 14.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 199.700 1.120 202.940 ;
  LAYER metal4 ;
  RECT 0.000 199.700 1.120 202.940 ;
  LAYER metal3 ;
  RECT 0.000 199.700 1.120 202.940 ;
  LAYER metal2 ;
  RECT 0.000 199.700 1.120 202.940 ;
  LAYER metal1 ;
  RECT 0.000 199.700 1.120 202.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 191.860 1.120 195.100 ;
  LAYER metal4 ;
  RECT 0.000 191.860 1.120 195.100 ;
  LAYER metal3 ;
  RECT 0.000 191.860 1.120 195.100 ;
  LAYER metal2 ;
  RECT 0.000 191.860 1.120 195.100 ;
  LAYER metal1 ;
  RECT 0.000 191.860 1.120 195.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 184.020 1.120 187.260 ;
  LAYER metal4 ;
  RECT 0.000 184.020 1.120 187.260 ;
  LAYER metal3 ;
  RECT 0.000 184.020 1.120 187.260 ;
  LAYER metal2 ;
  RECT 0.000 184.020 1.120 187.260 ;
  LAYER metal1 ;
  RECT 0.000 184.020 1.120 187.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 176.180 1.120 179.420 ;
  LAYER metal4 ;
  RECT 0.000 176.180 1.120 179.420 ;
  LAYER metal3 ;
  RECT 0.000 176.180 1.120 179.420 ;
  LAYER metal2 ;
  RECT 0.000 176.180 1.120 179.420 ;
  LAYER metal1 ;
  RECT 0.000 176.180 1.120 179.420 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 168.340 1.120 171.580 ;
  LAYER metal4 ;
  RECT 0.000 168.340 1.120 171.580 ;
  LAYER metal3 ;
  RECT 0.000 168.340 1.120 171.580 ;
  LAYER metal2 ;
  RECT 0.000 168.340 1.120 171.580 ;
  LAYER metal1 ;
  RECT 0.000 168.340 1.120 171.580 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 129.140 1.120 132.380 ;
  LAYER metal4 ;
  RECT 0.000 129.140 1.120 132.380 ;
  LAYER metal3 ;
  RECT 0.000 129.140 1.120 132.380 ;
  LAYER metal2 ;
  RECT 0.000 129.140 1.120 132.380 ;
  LAYER metal1 ;
  RECT 0.000 129.140 1.120 132.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 121.300 1.120 124.540 ;
  LAYER metal4 ;
  RECT 0.000 121.300 1.120 124.540 ;
  LAYER metal3 ;
  RECT 0.000 121.300 1.120 124.540 ;
  LAYER metal2 ;
  RECT 0.000 121.300 1.120 124.540 ;
  LAYER metal1 ;
  RECT 0.000 121.300 1.120 124.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 113.460 1.120 116.700 ;
  LAYER metal4 ;
  RECT 0.000 113.460 1.120 116.700 ;
  LAYER metal3 ;
  RECT 0.000 113.460 1.120 116.700 ;
  LAYER metal2 ;
  RECT 0.000 113.460 1.120 116.700 ;
  LAYER metal1 ;
  RECT 0.000 113.460 1.120 116.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 105.620 1.120 108.860 ;
  LAYER metal4 ;
  RECT 0.000 105.620 1.120 108.860 ;
  LAYER metal3 ;
  RECT 0.000 105.620 1.120 108.860 ;
  LAYER metal2 ;
  RECT 0.000 105.620 1.120 108.860 ;
  LAYER metal1 ;
  RECT 0.000 105.620 1.120 108.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 97.780 1.120 101.020 ;
  LAYER metal4 ;
  RECT 0.000 97.780 1.120 101.020 ;
  LAYER metal3 ;
  RECT 0.000 97.780 1.120 101.020 ;
  LAYER metal2 ;
  RECT 0.000 97.780 1.120 101.020 ;
  LAYER metal1 ;
  RECT 0.000 97.780 1.120 101.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 89.940 1.120 93.180 ;
  LAYER metal4 ;
  RECT 0.000 89.940 1.120 93.180 ;
  LAYER metal3 ;
  RECT 0.000 89.940 1.120 93.180 ;
  LAYER metal2 ;
  RECT 0.000 89.940 1.120 93.180 ;
  LAYER metal1 ;
  RECT 0.000 89.940 1.120 93.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 50.740 1.120 53.980 ;
  LAYER metal4 ;
  RECT 0.000 50.740 1.120 53.980 ;
  LAYER metal3 ;
  RECT 0.000 50.740 1.120 53.980 ;
  LAYER metal2 ;
  RECT 0.000 50.740 1.120 53.980 ;
  LAYER metal1 ;
  RECT 0.000 50.740 1.120 53.980 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 42.900 1.120 46.140 ;
  LAYER metal4 ;
  RECT 0.000 42.900 1.120 46.140 ;
  LAYER metal3 ;
  RECT 0.000 42.900 1.120 46.140 ;
  LAYER metal2 ;
  RECT 0.000 42.900 1.120 46.140 ;
  LAYER metal1 ;
  RECT 0.000 42.900 1.120 46.140 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 35.060 1.120 38.300 ;
  LAYER metal4 ;
  RECT 0.000 35.060 1.120 38.300 ;
  LAYER metal3 ;
  RECT 0.000 35.060 1.120 38.300 ;
  LAYER metal2 ;
  RECT 0.000 35.060 1.120 38.300 ;
  LAYER metal1 ;
  RECT 0.000 35.060 1.120 38.300 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 27.220 1.120 30.460 ;
  LAYER metal4 ;
  RECT 0.000 27.220 1.120 30.460 ;
  LAYER metal3 ;
  RECT 0.000 27.220 1.120 30.460 ;
  LAYER metal2 ;
  RECT 0.000 27.220 1.120 30.460 ;
  LAYER metal1 ;
  RECT 0.000 27.220 1.120 30.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 19.380 1.120 22.620 ;
  LAYER metal4 ;
  RECT 0.000 19.380 1.120 22.620 ;
  LAYER metal3 ;
  RECT 0.000 19.380 1.120 22.620 ;
  LAYER metal2 ;
  RECT 0.000 19.380 1.120 22.620 ;
  LAYER metal1 ;
  RECT 0.000 19.380 1.120 22.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 11.540 1.120 14.780 ;
  LAYER metal4 ;
  RECT 0.000 11.540 1.120 14.780 ;
  LAYER metal3 ;
  RECT 0.000 11.540 1.120 14.780 ;
  LAYER metal2 ;
  RECT 0.000 11.540 1.120 14.780 ;
  LAYER metal1 ;
  RECT 0.000 11.540 1.120 14.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3555.480 208.880 3559.020 210.000 ;
  LAYER metal4 ;
  RECT 3555.480 208.880 3559.020 210.000 ;
  LAYER metal3 ;
  RECT 3555.480 208.880 3559.020 210.000 ;
  LAYER metal2 ;
  RECT 3555.480 208.880 3559.020 210.000 ;
  LAYER metal1 ;
  RECT 3555.480 208.880 3559.020 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3541.840 208.880 3545.380 210.000 ;
  LAYER metal4 ;
  RECT 3541.840 208.880 3545.380 210.000 ;
  LAYER metal3 ;
  RECT 3541.840 208.880 3545.380 210.000 ;
  LAYER metal2 ;
  RECT 3541.840 208.880 3545.380 210.000 ;
  LAYER metal1 ;
  RECT 3541.840 208.880 3545.380 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3528.820 208.880 3532.360 210.000 ;
  LAYER metal4 ;
  RECT 3528.820 208.880 3532.360 210.000 ;
  LAYER metal3 ;
  RECT 3528.820 208.880 3532.360 210.000 ;
  LAYER metal2 ;
  RECT 3528.820 208.880 3532.360 210.000 ;
  LAYER metal1 ;
  RECT 3528.820 208.880 3532.360 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3461.240 208.880 3464.780 210.000 ;
  LAYER metal4 ;
  RECT 3461.240 208.880 3464.780 210.000 ;
  LAYER metal3 ;
  RECT 3461.240 208.880 3464.780 210.000 ;
  LAYER metal2 ;
  RECT 3461.240 208.880 3464.780 210.000 ;
  LAYER metal1 ;
  RECT 3461.240 208.880 3464.780 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3447.600 208.880 3451.140 210.000 ;
  LAYER metal4 ;
  RECT 3447.600 208.880 3451.140 210.000 ;
  LAYER metal3 ;
  RECT 3447.600 208.880 3451.140 210.000 ;
  LAYER metal2 ;
  RECT 3447.600 208.880 3451.140 210.000 ;
  LAYER metal1 ;
  RECT 3447.600 208.880 3451.140 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3434.580 208.880 3438.120 210.000 ;
  LAYER metal4 ;
  RECT 3434.580 208.880 3438.120 210.000 ;
  LAYER metal3 ;
  RECT 3434.580 208.880 3438.120 210.000 ;
  LAYER metal2 ;
  RECT 3434.580 208.880 3438.120 210.000 ;
  LAYER metal1 ;
  RECT 3434.580 208.880 3438.120 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3420.940 208.880 3424.480 210.000 ;
  LAYER metal4 ;
  RECT 3420.940 208.880 3424.480 210.000 ;
  LAYER metal3 ;
  RECT 3420.940 208.880 3424.480 210.000 ;
  LAYER metal2 ;
  RECT 3420.940 208.880 3424.480 210.000 ;
  LAYER metal1 ;
  RECT 3420.940 208.880 3424.480 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3407.300 208.880 3410.840 210.000 ;
  LAYER metal4 ;
  RECT 3407.300 208.880 3410.840 210.000 ;
  LAYER metal3 ;
  RECT 3407.300 208.880 3410.840 210.000 ;
  LAYER metal2 ;
  RECT 3407.300 208.880 3410.840 210.000 ;
  LAYER metal1 ;
  RECT 3407.300 208.880 3410.840 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3394.280 208.880 3397.820 210.000 ;
  LAYER metal4 ;
  RECT 3394.280 208.880 3397.820 210.000 ;
  LAYER metal3 ;
  RECT 3394.280 208.880 3397.820 210.000 ;
  LAYER metal2 ;
  RECT 3394.280 208.880 3397.820 210.000 ;
  LAYER metal1 ;
  RECT 3394.280 208.880 3397.820 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3326.700 208.880 3330.240 210.000 ;
  LAYER metal4 ;
  RECT 3326.700 208.880 3330.240 210.000 ;
  LAYER metal3 ;
  RECT 3326.700 208.880 3330.240 210.000 ;
  LAYER metal2 ;
  RECT 3326.700 208.880 3330.240 210.000 ;
  LAYER metal1 ;
  RECT 3326.700 208.880 3330.240 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3313.680 208.880 3317.220 210.000 ;
  LAYER metal4 ;
  RECT 3313.680 208.880 3317.220 210.000 ;
  LAYER metal3 ;
  RECT 3313.680 208.880 3317.220 210.000 ;
  LAYER metal2 ;
  RECT 3313.680 208.880 3317.220 210.000 ;
  LAYER metal1 ;
  RECT 3313.680 208.880 3317.220 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3300.040 208.880 3303.580 210.000 ;
  LAYER metal4 ;
  RECT 3300.040 208.880 3303.580 210.000 ;
  LAYER metal3 ;
  RECT 3300.040 208.880 3303.580 210.000 ;
  LAYER metal2 ;
  RECT 3300.040 208.880 3303.580 210.000 ;
  LAYER metal1 ;
  RECT 3300.040 208.880 3303.580 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3286.400 208.880 3289.940 210.000 ;
  LAYER metal4 ;
  RECT 3286.400 208.880 3289.940 210.000 ;
  LAYER metal3 ;
  RECT 3286.400 208.880 3289.940 210.000 ;
  LAYER metal2 ;
  RECT 3286.400 208.880 3289.940 210.000 ;
  LAYER metal1 ;
  RECT 3286.400 208.880 3289.940 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3273.380 208.880 3276.920 210.000 ;
  LAYER metal4 ;
  RECT 3273.380 208.880 3276.920 210.000 ;
  LAYER metal3 ;
  RECT 3273.380 208.880 3276.920 210.000 ;
  LAYER metal2 ;
  RECT 3273.380 208.880 3276.920 210.000 ;
  LAYER metal1 ;
  RECT 3273.380 208.880 3276.920 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3259.740 208.880 3263.280 210.000 ;
  LAYER metal4 ;
  RECT 3259.740 208.880 3263.280 210.000 ;
  LAYER metal3 ;
  RECT 3259.740 208.880 3263.280 210.000 ;
  LAYER metal2 ;
  RECT 3259.740 208.880 3263.280 210.000 ;
  LAYER metal1 ;
  RECT 3259.740 208.880 3263.280 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3192.780 208.880 3196.320 210.000 ;
  LAYER metal4 ;
  RECT 3192.780 208.880 3196.320 210.000 ;
  LAYER metal3 ;
  RECT 3192.780 208.880 3196.320 210.000 ;
  LAYER metal2 ;
  RECT 3192.780 208.880 3196.320 210.000 ;
  LAYER metal1 ;
  RECT 3192.780 208.880 3196.320 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3179.140 208.880 3182.680 210.000 ;
  LAYER metal4 ;
  RECT 3179.140 208.880 3182.680 210.000 ;
  LAYER metal3 ;
  RECT 3179.140 208.880 3182.680 210.000 ;
  LAYER metal2 ;
  RECT 3179.140 208.880 3182.680 210.000 ;
  LAYER metal1 ;
  RECT 3179.140 208.880 3182.680 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3165.500 208.880 3169.040 210.000 ;
  LAYER metal4 ;
  RECT 3165.500 208.880 3169.040 210.000 ;
  LAYER metal3 ;
  RECT 3165.500 208.880 3169.040 210.000 ;
  LAYER metal2 ;
  RECT 3165.500 208.880 3169.040 210.000 ;
  LAYER metal1 ;
  RECT 3165.500 208.880 3169.040 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3152.480 208.880 3156.020 210.000 ;
  LAYER metal4 ;
  RECT 3152.480 208.880 3156.020 210.000 ;
  LAYER metal3 ;
  RECT 3152.480 208.880 3156.020 210.000 ;
  LAYER metal2 ;
  RECT 3152.480 208.880 3156.020 210.000 ;
  LAYER metal1 ;
  RECT 3152.480 208.880 3156.020 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3138.840 208.880 3142.380 210.000 ;
  LAYER metal4 ;
  RECT 3138.840 208.880 3142.380 210.000 ;
  LAYER metal3 ;
  RECT 3138.840 208.880 3142.380 210.000 ;
  LAYER metal2 ;
  RECT 3138.840 208.880 3142.380 210.000 ;
  LAYER metal1 ;
  RECT 3138.840 208.880 3142.380 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3125.200 208.880 3128.740 210.000 ;
  LAYER metal4 ;
  RECT 3125.200 208.880 3128.740 210.000 ;
  LAYER metal3 ;
  RECT 3125.200 208.880 3128.740 210.000 ;
  LAYER metal2 ;
  RECT 3125.200 208.880 3128.740 210.000 ;
  LAYER metal1 ;
  RECT 3125.200 208.880 3128.740 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3058.240 208.880 3061.780 210.000 ;
  LAYER metal4 ;
  RECT 3058.240 208.880 3061.780 210.000 ;
  LAYER metal3 ;
  RECT 3058.240 208.880 3061.780 210.000 ;
  LAYER metal2 ;
  RECT 3058.240 208.880 3061.780 210.000 ;
  LAYER metal1 ;
  RECT 3058.240 208.880 3061.780 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3044.600 208.880 3048.140 210.000 ;
  LAYER metal4 ;
  RECT 3044.600 208.880 3048.140 210.000 ;
  LAYER metal3 ;
  RECT 3044.600 208.880 3048.140 210.000 ;
  LAYER metal2 ;
  RECT 3044.600 208.880 3048.140 210.000 ;
  LAYER metal1 ;
  RECT 3044.600 208.880 3048.140 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3030.960 208.880 3034.500 210.000 ;
  LAYER metal4 ;
  RECT 3030.960 208.880 3034.500 210.000 ;
  LAYER metal3 ;
  RECT 3030.960 208.880 3034.500 210.000 ;
  LAYER metal2 ;
  RECT 3030.960 208.880 3034.500 210.000 ;
  LAYER metal1 ;
  RECT 3030.960 208.880 3034.500 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3017.940 208.880 3021.480 210.000 ;
  LAYER metal4 ;
  RECT 3017.940 208.880 3021.480 210.000 ;
  LAYER metal3 ;
  RECT 3017.940 208.880 3021.480 210.000 ;
  LAYER metal2 ;
  RECT 3017.940 208.880 3021.480 210.000 ;
  LAYER metal1 ;
  RECT 3017.940 208.880 3021.480 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3004.300 208.880 3007.840 210.000 ;
  LAYER metal4 ;
  RECT 3004.300 208.880 3007.840 210.000 ;
  LAYER metal3 ;
  RECT 3004.300 208.880 3007.840 210.000 ;
  LAYER metal2 ;
  RECT 3004.300 208.880 3007.840 210.000 ;
  LAYER metal1 ;
  RECT 3004.300 208.880 3007.840 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2990.660 208.880 2994.200 210.000 ;
  LAYER metal4 ;
  RECT 2990.660 208.880 2994.200 210.000 ;
  LAYER metal3 ;
  RECT 2990.660 208.880 2994.200 210.000 ;
  LAYER metal2 ;
  RECT 2990.660 208.880 2994.200 210.000 ;
  LAYER metal1 ;
  RECT 2990.660 208.880 2994.200 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2923.700 208.880 2927.240 210.000 ;
  LAYER metal4 ;
  RECT 2923.700 208.880 2927.240 210.000 ;
  LAYER metal3 ;
  RECT 2923.700 208.880 2927.240 210.000 ;
  LAYER metal2 ;
  RECT 2923.700 208.880 2927.240 210.000 ;
  LAYER metal1 ;
  RECT 2923.700 208.880 2927.240 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2910.060 208.880 2913.600 210.000 ;
  LAYER metal4 ;
  RECT 2910.060 208.880 2913.600 210.000 ;
  LAYER metal3 ;
  RECT 2910.060 208.880 2913.600 210.000 ;
  LAYER metal2 ;
  RECT 2910.060 208.880 2913.600 210.000 ;
  LAYER metal1 ;
  RECT 2910.060 208.880 2913.600 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2897.040 208.880 2900.580 210.000 ;
  LAYER metal4 ;
  RECT 2897.040 208.880 2900.580 210.000 ;
  LAYER metal3 ;
  RECT 2897.040 208.880 2900.580 210.000 ;
  LAYER metal2 ;
  RECT 2897.040 208.880 2900.580 210.000 ;
  LAYER metal1 ;
  RECT 2897.040 208.880 2900.580 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2883.400 208.880 2886.940 210.000 ;
  LAYER metal4 ;
  RECT 2883.400 208.880 2886.940 210.000 ;
  LAYER metal3 ;
  RECT 2883.400 208.880 2886.940 210.000 ;
  LAYER metal2 ;
  RECT 2883.400 208.880 2886.940 210.000 ;
  LAYER metal1 ;
  RECT 2883.400 208.880 2886.940 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2869.760 208.880 2873.300 210.000 ;
  LAYER metal4 ;
  RECT 2869.760 208.880 2873.300 210.000 ;
  LAYER metal3 ;
  RECT 2869.760 208.880 2873.300 210.000 ;
  LAYER metal2 ;
  RECT 2869.760 208.880 2873.300 210.000 ;
  LAYER metal1 ;
  RECT 2869.760 208.880 2873.300 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2856.740 208.880 2860.280 210.000 ;
  LAYER metal4 ;
  RECT 2856.740 208.880 2860.280 210.000 ;
  LAYER metal3 ;
  RECT 2856.740 208.880 2860.280 210.000 ;
  LAYER metal2 ;
  RECT 2856.740 208.880 2860.280 210.000 ;
  LAYER metal1 ;
  RECT 2856.740 208.880 2860.280 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2789.160 208.880 2792.700 210.000 ;
  LAYER metal4 ;
  RECT 2789.160 208.880 2792.700 210.000 ;
  LAYER metal3 ;
  RECT 2789.160 208.880 2792.700 210.000 ;
  LAYER metal2 ;
  RECT 2789.160 208.880 2792.700 210.000 ;
  LAYER metal1 ;
  RECT 2789.160 208.880 2792.700 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2776.140 208.880 2779.680 210.000 ;
  LAYER metal4 ;
  RECT 2776.140 208.880 2779.680 210.000 ;
  LAYER metal3 ;
  RECT 2776.140 208.880 2779.680 210.000 ;
  LAYER metal2 ;
  RECT 2776.140 208.880 2779.680 210.000 ;
  LAYER metal1 ;
  RECT 2776.140 208.880 2779.680 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2762.500 208.880 2766.040 210.000 ;
  LAYER metal4 ;
  RECT 2762.500 208.880 2766.040 210.000 ;
  LAYER metal3 ;
  RECT 2762.500 208.880 2766.040 210.000 ;
  LAYER metal2 ;
  RECT 2762.500 208.880 2766.040 210.000 ;
  LAYER metal1 ;
  RECT 2762.500 208.880 2766.040 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2748.860 208.880 2752.400 210.000 ;
  LAYER metal4 ;
  RECT 2748.860 208.880 2752.400 210.000 ;
  LAYER metal3 ;
  RECT 2748.860 208.880 2752.400 210.000 ;
  LAYER metal2 ;
  RECT 2748.860 208.880 2752.400 210.000 ;
  LAYER metal1 ;
  RECT 2748.860 208.880 2752.400 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2735.840 208.880 2739.380 210.000 ;
  LAYER metal4 ;
  RECT 2735.840 208.880 2739.380 210.000 ;
  LAYER metal3 ;
  RECT 2735.840 208.880 2739.380 210.000 ;
  LAYER metal2 ;
  RECT 2735.840 208.880 2739.380 210.000 ;
  LAYER metal1 ;
  RECT 2735.840 208.880 2739.380 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2722.200 208.880 2725.740 210.000 ;
  LAYER metal4 ;
  RECT 2722.200 208.880 2725.740 210.000 ;
  LAYER metal3 ;
  RECT 2722.200 208.880 2725.740 210.000 ;
  LAYER metal2 ;
  RECT 2722.200 208.880 2725.740 210.000 ;
  LAYER metal1 ;
  RECT 2722.200 208.880 2725.740 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2655.240 208.880 2658.780 210.000 ;
  LAYER metal4 ;
  RECT 2655.240 208.880 2658.780 210.000 ;
  LAYER metal3 ;
  RECT 2655.240 208.880 2658.780 210.000 ;
  LAYER metal2 ;
  RECT 2655.240 208.880 2658.780 210.000 ;
  LAYER metal1 ;
  RECT 2655.240 208.880 2658.780 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2641.600 208.880 2645.140 210.000 ;
  LAYER metal4 ;
  RECT 2641.600 208.880 2645.140 210.000 ;
  LAYER metal3 ;
  RECT 2641.600 208.880 2645.140 210.000 ;
  LAYER metal2 ;
  RECT 2641.600 208.880 2645.140 210.000 ;
  LAYER metal1 ;
  RECT 2641.600 208.880 2645.140 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2627.960 208.880 2631.500 210.000 ;
  LAYER metal4 ;
  RECT 2627.960 208.880 2631.500 210.000 ;
  LAYER metal3 ;
  RECT 2627.960 208.880 2631.500 210.000 ;
  LAYER metal2 ;
  RECT 2627.960 208.880 2631.500 210.000 ;
  LAYER metal1 ;
  RECT 2627.960 208.880 2631.500 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2614.320 208.880 2617.860 210.000 ;
  LAYER metal4 ;
  RECT 2614.320 208.880 2617.860 210.000 ;
  LAYER metal3 ;
  RECT 2614.320 208.880 2617.860 210.000 ;
  LAYER metal2 ;
  RECT 2614.320 208.880 2617.860 210.000 ;
  LAYER metal1 ;
  RECT 2614.320 208.880 2617.860 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2601.300 208.880 2604.840 210.000 ;
  LAYER metal4 ;
  RECT 2601.300 208.880 2604.840 210.000 ;
  LAYER metal3 ;
  RECT 2601.300 208.880 2604.840 210.000 ;
  LAYER metal2 ;
  RECT 2601.300 208.880 2604.840 210.000 ;
  LAYER metal1 ;
  RECT 2601.300 208.880 2604.840 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2587.660 208.880 2591.200 210.000 ;
  LAYER metal4 ;
  RECT 2587.660 208.880 2591.200 210.000 ;
  LAYER metal3 ;
  RECT 2587.660 208.880 2591.200 210.000 ;
  LAYER metal2 ;
  RECT 2587.660 208.880 2591.200 210.000 ;
  LAYER metal1 ;
  RECT 2587.660 208.880 2591.200 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2520.700 208.880 2524.240 210.000 ;
  LAYER metal4 ;
  RECT 2520.700 208.880 2524.240 210.000 ;
  LAYER metal3 ;
  RECT 2520.700 208.880 2524.240 210.000 ;
  LAYER metal2 ;
  RECT 2520.700 208.880 2524.240 210.000 ;
  LAYER metal1 ;
  RECT 2520.700 208.880 2524.240 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2507.060 208.880 2510.600 210.000 ;
  LAYER metal4 ;
  RECT 2507.060 208.880 2510.600 210.000 ;
  LAYER metal3 ;
  RECT 2507.060 208.880 2510.600 210.000 ;
  LAYER metal2 ;
  RECT 2507.060 208.880 2510.600 210.000 ;
  LAYER metal1 ;
  RECT 2507.060 208.880 2510.600 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2493.420 208.880 2496.960 210.000 ;
  LAYER metal4 ;
  RECT 2493.420 208.880 2496.960 210.000 ;
  LAYER metal3 ;
  RECT 2493.420 208.880 2496.960 210.000 ;
  LAYER metal2 ;
  RECT 2493.420 208.880 2496.960 210.000 ;
  LAYER metal1 ;
  RECT 2493.420 208.880 2496.960 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2480.400 208.880 2483.940 210.000 ;
  LAYER metal4 ;
  RECT 2480.400 208.880 2483.940 210.000 ;
  LAYER metal3 ;
  RECT 2480.400 208.880 2483.940 210.000 ;
  LAYER metal2 ;
  RECT 2480.400 208.880 2483.940 210.000 ;
  LAYER metal1 ;
  RECT 2480.400 208.880 2483.940 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2466.760 208.880 2470.300 210.000 ;
  LAYER metal4 ;
  RECT 2466.760 208.880 2470.300 210.000 ;
  LAYER metal3 ;
  RECT 2466.760 208.880 2470.300 210.000 ;
  LAYER metal2 ;
  RECT 2466.760 208.880 2470.300 210.000 ;
  LAYER metal1 ;
  RECT 2466.760 208.880 2470.300 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2453.120 208.880 2456.660 210.000 ;
  LAYER metal4 ;
  RECT 2453.120 208.880 2456.660 210.000 ;
  LAYER metal3 ;
  RECT 2453.120 208.880 2456.660 210.000 ;
  LAYER metal2 ;
  RECT 2453.120 208.880 2456.660 210.000 ;
  LAYER metal1 ;
  RECT 2453.120 208.880 2456.660 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2386.160 208.880 2389.700 210.000 ;
  LAYER metal4 ;
  RECT 2386.160 208.880 2389.700 210.000 ;
  LAYER metal3 ;
  RECT 2386.160 208.880 2389.700 210.000 ;
  LAYER metal2 ;
  RECT 2386.160 208.880 2389.700 210.000 ;
  LAYER metal1 ;
  RECT 2386.160 208.880 2389.700 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2372.520 208.880 2376.060 210.000 ;
  LAYER metal4 ;
  RECT 2372.520 208.880 2376.060 210.000 ;
  LAYER metal3 ;
  RECT 2372.520 208.880 2376.060 210.000 ;
  LAYER metal2 ;
  RECT 2372.520 208.880 2376.060 210.000 ;
  LAYER metal1 ;
  RECT 2372.520 208.880 2376.060 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2359.500 208.880 2363.040 210.000 ;
  LAYER metal4 ;
  RECT 2359.500 208.880 2363.040 210.000 ;
  LAYER metal3 ;
  RECT 2359.500 208.880 2363.040 210.000 ;
  LAYER metal2 ;
  RECT 2359.500 208.880 2363.040 210.000 ;
  LAYER metal1 ;
  RECT 2359.500 208.880 2363.040 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2345.860 208.880 2349.400 210.000 ;
  LAYER metal4 ;
  RECT 2345.860 208.880 2349.400 210.000 ;
  LAYER metal3 ;
  RECT 2345.860 208.880 2349.400 210.000 ;
  LAYER metal2 ;
  RECT 2345.860 208.880 2349.400 210.000 ;
  LAYER metal1 ;
  RECT 2345.860 208.880 2349.400 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2332.220 208.880 2335.760 210.000 ;
  LAYER metal4 ;
  RECT 2332.220 208.880 2335.760 210.000 ;
  LAYER metal3 ;
  RECT 2332.220 208.880 2335.760 210.000 ;
  LAYER metal2 ;
  RECT 2332.220 208.880 2335.760 210.000 ;
  LAYER metal1 ;
  RECT 2332.220 208.880 2335.760 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2319.200 208.880 2322.740 210.000 ;
  LAYER metal4 ;
  RECT 2319.200 208.880 2322.740 210.000 ;
  LAYER metal3 ;
  RECT 2319.200 208.880 2322.740 210.000 ;
  LAYER metal2 ;
  RECT 2319.200 208.880 2322.740 210.000 ;
  LAYER metal1 ;
  RECT 2319.200 208.880 2322.740 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2251.620 208.880 2255.160 210.000 ;
  LAYER metal4 ;
  RECT 2251.620 208.880 2255.160 210.000 ;
  LAYER metal3 ;
  RECT 2251.620 208.880 2255.160 210.000 ;
  LAYER metal2 ;
  RECT 2251.620 208.880 2255.160 210.000 ;
  LAYER metal1 ;
  RECT 2251.620 208.880 2255.160 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2238.600 208.880 2242.140 210.000 ;
  LAYER metal4 ;
  RECT 2238.600 208.880 2242.140 210.000 ;
  LAYER metal3 ;
  RECT 2238.600 208.880 2242.140 210.000 ;
  LAYER metal2 ;
  RECT 2238.600 208.880 2242.140 210.000 ;
  LAYER metal1 ;
  RECT 2238.600 208.880 2242.140 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2224.960 208.880 2228.500 210.000 ;
  LAYER metal4 ;
  RECT 2224.960 208.880 2228.500 210.000 ;
  LAYER metal3 ;
  RECT 2224.960 208.880 2228.500 210.000 ;
  LAYER metal2 ;
  RECT 2224.960 208.880 2228.500 210.000 ;
  LAYER metal1 ;
  RECT 2224.960 208.880 2228.500 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2211.320 208.880 2214.860 210.000 ;
  LAYER metal4 ;
  RECT 2211.320 208.880 2214.860 210.000 ;
  LAYER metal3 ;
  RECT 2211.320 208.880 2214.860 210.000 ;
  LAYER metal2 ;
  RECT 2211.320 208.880 2214.860 210.000 ;
  LAYER metal1 ;
  RECT 2211.320 208.880 2214.860 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2197.680 208.880 2201.220 210.000 ;
  LAYER metal4 ;
  RECT 2197.680 208.880 2201.220 210.000 ;
  LAYER metal3 ;
  RECT 2197.680 208.880 2201.220 210.000 ;
  LAYER metal2 ;
  RECT 2197.680 208.880 2201.220 210.000 ;
  LAYER metal1 ;
  RECT 2197.680 208.880 2201.220 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2184.660 208.880 2188.200 210.000 ;
  LAYER metal4 ;
  RECT 2184.660 208.880 2188.200 210.000 ;
  LAYER metal3 ;
  RECT 2184.660 208.880 2188.200 210.000 ;
  LAYER metal2 ;
  RECT 2184.660 208.880 2188.200 210.000 ;
  LAYER metal1 ;
  RECT 2184.660 208.880 2188.200 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2117.080 208.880 2120.620 210.000 ;
  LAYER metal4 ;
  RECT 2117.080 208.880 2120.620 210.000 ;
  LAYER metal3 ;
  RECT 2117.080 208.880 2120.620 210.000 ;
  LAYER metal2 ;
  RECT 2117.080 208.880 2120.620 210.000 ;
  LAYER metal1 ;
  RECT 2117.080 208.880 2120.620 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2104.060 208.880 2107.600 210.000 ;
  LAYER metal4 ;
  RECT 2104.060 208.880 2107.600 210.000 ;
  LAYER metal3 ;
  RECT 2104.060 208.880 2107.600 210.000 ;
  LAYER metal2 ;
  RECT 2104.060 208.880 2107.600 210.000 ;
  LAYER metal1 ;
  RECT 2104.060 208.880 2107.600 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2090.420 208.880 2093.960 210.000 ;
  LAYER metal4 ;
  RECT 2090.420 208.880 2093.960 210.000 ;
  LAYER metal3 ;
  RECT 2090.420 208.880 2093.960 210.000 ;
  LAYER metal2 ;
  RECT 2090.420 208.880 2093.960 210.000 ;
  LAYER metal1 ;
  RECT 2090.420 208.880 2093.960 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2076.780 208.880 2080.320 210.000 ;
  LAYER metal4 ;
  RECT 2076.780 208.880 2080.320 210.000 ;
  LAYER metal3 ;
  RECT 2076.780 208.880 2080.320 210.000 ;
  LAYER metal2 ;
  RECT 2076.780 208.880 2080.320 210.000 ;
  LAYER metal1 ;
  RECT 2076.780 208.880 2080.320 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2063.760 208.880 2067.300 210.000 ;
  LAYER metal4 ;
  RECT 2063.760 208.880 2067.300 210.000 ;
  LAYER metal3 ;
  RECT 2063.760 208.880 2067.300 210.000 ;
  LAYER metal2 ;
  RECT 2063.760 208.880 2067.300 210.000 ;
  LAYER metal1 ;
  RECT 2063.760 208.880 2067.300 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2050.120 208.880 2053.660 210.000 ;
  LAYER metal4 ;
  RECT 2050.120 208.880 2053.660 210.000 ;
  LAYER metal3 ;
  RECT 2050.120 208.880 2053.660 210.000 ;
  LAYER metal2 ;
  RECT 2050.120 208.880 2053.660 210.000 ;
  LAYER metal1 ;
  RECT 2050.120 208.880 2053.660 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1983.160 208.880 1986.700 210.000 ;
  LAYER metal4 ;
  RECT 1983.160 208.880 1986.700 210.000 ;
  LAYER metal3 ;
  RECT 1983.160 208.880 1986.700 210.000 ;
  LAYER metal2 ;
  RECT 1983.160 208.880 1986.700 210.000 ;
  LAYER metal1 ;
  RECT 1983.160 208.880 1986.700 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1969.520 208.880 1973.060 210.000 ;
  LAYER metal4 ;
  RECT 1969.520 208.880 1973.060 210.000 ;
  LAYER metal3 ;
  RECT 1969.520 208.880 1973.060 210.000 ;
  LAYER metal2 ;
  RECT 1969.520 208.880 1973.060 210.000 ;
  LAYER metal1 ;
  RECT 1969.520 208.880 1973.060 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1955.880 208.880 1959.420 210.000 ;
  LAYER metal4 ;
  RECT 1955.880 208.880 1959.420 210.000 ;
  LAYER metal3 ;
  RECT 1955.880 208.880 1959.420 210.000 ;
  LAYER metal2 ;
  RECT 1955.880 208.880 1959.420 210.000 ;
  LAYER metal1 ;
  RECT 1955.880 208.880 1959.420 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1942.860 208.880 1946.400 210.000 ;
  LAYER metal4 ;
  RECT 1942.860 208.880 1946.400 210.000 ;
  LAYER metal3 ;
  RECT 1942.860 208.880 1946.400 210.000 ;
  LAYER metal2 ;
  RECT 1942.860 208.880 1946.400 210.000 ;
  LAYER metal1 ;
  RECT 1942.860 208.880 1946.400 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1929.220 208.880 1932.760 210.000 ;
  LAYER metal4 ;
  RECT 1929.220 208.880 1932.760 210.000 ;
  LAYER metal3 ;
  RECT 1929.220 208.880 1932.760 210.000 ;
  LAYER metal2 ;
  RECT 1929.220 208.880 1932.760 210.000 ;
  LAYER metal1 ;
  RECT 1929.220 208.880 1932.760 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1915.580 208.880 1919.120 210.000 ;
  LAYER metal4 ;
  RECT 1915.580 208.880 1919.120 210.000 ;
  LAYER metal3 ;
  RECT 1915.580 208.880 1919.120 210.000 ;
  LAYER metal2 ;
  RECT 1915.580 208.880 1919.120 210.000 ;
  LAYER metal1 ;
  RECT 1915.580 208.880 1919.120 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1848.620 208.880 1852.160 210.000 ;
  LAYER metal4 ;
  RECT 1848.620 208.880 1852.160 210.000 ;
  LAYER metal3 ;
  RECT 1848.620 208.880 1852.160 210.000 ;
  LAYER metal2 ;
  RECT 1848.620 208.880 1852.160 210.000 ;
  LAYER metal1 ;
  RECT 1848.620 208.880 1852.160 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1834.980 208.880 1838.520 210.000 ;
  LAYER metal4 ;
  RECT 1834.980 208.880 1838.520 210.000 ;
  LAYER metal3 ;
  RECT 1834.980 208.880 1838.520 210.000 ;
  LAYER metal2 ;
  RECT 1834.980 208.880 1838.520 210.000 ;
  LAYER metal1 ;
  RECT 1834.980 208.880 1838.520 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1826.300 208.880 1829.840 210.000 ;
  LAYER metal4 ;
  RECT 1826.300 208.880 1829.840 210.000 ;
  LAYER metal3 ;
  RECT 1826.300 208.880 1829.840 210.000 ;
  LAYER metal2 ;
  RECT 1826.300 208.880 1829.840 210.000 ;
  LAYER metal1 ;
  RECT 1826.300 208.880 1829.840 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1817.620 208.880 1821.160 210.000 ;
  LAYER metal4 ;
  RECT 1817.620 208.880 1821.160 210.000 ;
  LAYER metal3 ;
  RECT 1817.620 208.880 1821.160 210.000 ;
  LAYER metal2 ;
  RECT 1817.620 208.880 1821.160 210.000 ;
  LAYER metal1 ;
  RECT 1817.620 208.880 1821.160 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1803.980 208.880 1807.520 210.000 ;
  LAYER metal4 ;
  RECT 1803.980 208.880 1807.520 210.000 ;
  LAYER metal3 ;
  RECT 1803.980 208.880 1807.520 210.000 ;
  LAYER metal2 ;
  RECT 1803.980 208.880 1807.520 210.000 ;
  LAYER metal1 ;
  RECT 1803.980 208.880 1807.520 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1758.720 208.880 1762.260 210.000 ;
  LAYER metal4 ;
  RECT 1758.720 208.880 1762.260 210.000 ;
  LAYER metal3 ;
  RECT 1758.720 208.880 1762.260 210.000 ;
  LAYER metal2 ;
  RECT 1758.720 208.880 1762.260 210.000 ;
  LAYER metal1 ;
  RECT 1758.720 208.880 1762.260 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1694.860 208.880 1698.400 210.000 ;
  LAYER metal4 ;
  RECT 1694.860 208.880 1698.400 210.000 ;
  LAYER metal3 ;
  RECT 1694.860 208.880 1698.400 210.000 ;
  LAYER metal2 ;
  RECT 1694.860 208.880 1698.400 210.000 ;
  LAYER metal1 ;
  RECT 1694.860 208.880 1698.400 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1681.220 208.880 1684.760 210.000 ;
  LAYER metal4 ;
  RECT 1681.220 208.880 1684.760 210.000 ;
  LAYER metal3 ;
  RECT 1681.220 208.880 1684.760 210.000 ;
  LAYER metal2 ;
  RECT 1681.220 208.880 1684.760 210.000 ;
  LAYER metal1 ;
  RECT 1681.220 208.880 1684.760 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1668.200 208.880 1671.740 210.000 ;
  LAYER metal4 ;
  RECT 1668.200 208.880 1671.740 210.000 ;
  LAYER metal3 ;
  RECT 1668.200 208.880 1671.740 210.000 ;
  LAYER metal2 ;
  RECT 1668.200 208.880 1671.740 210.000 ;
  LAYER metal1 ;
  RECT 1668.200 208.880 1671.740 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1654.560 208.880 1658.100 210.000 ;
  LAYER metal4 ;
  RECT 1654.560 208.880 1658.100 210.000 ;
  LAYER metal3 ;
  RECT 1654.560 208.880 1658.100 210.000 ;
  LAYER metal2 ;
  RECT 1654.560 208.880 1658.100 210.000 ;
  LAYER metal1 ;
  RECT 1654.560 208.880 1658.100 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1640.920 208.880 1644.460 210.000 ;
  LAYER metal4 ;
  RECT 1640.920 208.880 1644.460 210.000 ;
  LAYER metal3 ;
  RECT 1640.920 208.880 1644.460 210.000 ;
  LAYER metal2 ;
  RECT 1640.920 208.880 1644.460 210.000 ;
  LAYER metal1 ;
  RECT 1640.920 208.880 1644.460 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1627.900 208.880 1631.440 210.000 ;
  LAYER metal4 ;
  RECT 1627.900 208.880 1631.440 210.000 ;
  LAYER metal3 ;
  RECT 1627.900 208.880 1631.440 210.000 ;
  LAYER metal2 ;
  RECT 1627.900 208.880 1631.440 210.000 ;
  LAYER metal1 ;
  RECT 1627.900 208.880 1631.440 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1560.320 208.880 1563.860 210.000 ;
  LAYER metal4 ;
  RECT 1560.320 208.880 1563.860 210.000 ;
  LAYER metal3 ;
  RECT 1560.320 208.880 1563.860 210.000 ;
  LAYER metal2 ;
  RECT 1560.320 208.880 1563.860 210.000 ;
  LAYER metal1 ;
  RECT 1560.320 208.880 1563.860 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1547.300 208.880 1550.840 210.000 ;
  LAYER metal4 ;
  RECT 1547.300 208.880 1550.840 210.000 ;
  LAYER metal3 ;
  RECT 1547.300 208.880 1550.840 210.000 ;
  LAYER metal2 ;
  RECT 1547.300 208.880 1550.840 210.000 ;
  LAYER metal1 ;
  RECT 1547.300 208.880 1550.840 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1533.660 208.880 1537.200 210.000 ;
  LAYER metal4 ;
  RECT 1533.660 208.880 1537.200 210.000 ;
  LAYER metal3 ;
  RECT 1533.660 208.880 1537.200 210.000 ;
  LAYER metal2 ;
  RECT 1533.660 208.880 1537.200 210.000 ;
  LAYER metal1 ;
  RECT 1533.660 208.880 1537.200 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1520.020 208.880 1523.560 210.000 ;
  LAYER metal4 ;
  RECT 1520.020 208.880 1523.560 210.000 ;
  LAYER metal3 ;
  RECT 1520.020 208.880 1523.560 210.000 ;
  LAYER metal2 ;
  RECT 1520.020 208.880 1523.560 210.000 ;
  LAYER metal1 ;
  RECT 1520.020 208.880 1523.560 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1507.000 208.880 1510.540 210.000 ;
  LAYER metal4 ;
  RECT 1507.000 208.880 1510.540 210.000 ;
  LAYER metal3 ;
  RECT 1507.000 208.880 1510.540 210.000 ;
  LAYER metal2 ;
  RECT 1507.000 208.880 1510.540 210.000 ;
  LAYER metal1 ;
  RECT 1507.000 208.880 1510.540 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1493.360 208.880 1496.900 210.000 ;
  LAYER metal4 ;
  RECT 1493.360 208.880 1496.900 210.000 ;
  LAYER metal3 ;
  RECT 1493.360 208.880 1496.900 210.000 ;
  LAYER metal2 ;
  RECT 1493.360 208.880 1496.900 210.000 ;
  LAYER metal1 ;
  RECT 1493.360 208.880 1496.900 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1426.400 208.880 1429.940 210.000 ;
  LAYER metal4 ;
  RECT 1426.400 208.880 1429.940 210.000 ;
  LAYER metal3 ;
  RECT 1426.400 208.880 1429.940 210.000 ;
  LAYER metal2 ;
  RECT 1426.400 208.880 1429.940 210.000 ;
  LAYER metal1 ;
  RECT 1426.400 208.880 1429.940 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1412.760 208.880 1416.300 210.000 ;
  LAYER metal4 ;
  RECT 1412.760 208.880 1416.300 210.000 ;
  LAYER metal3 ;
  RECT 1412.760 208.880 1416.300 210.000 ;
  LAYER metal2 ;
  RECT 1412.760 208.880 1416.300 210.000 ;
  LAYER metal1 ;
  RECT 1412.760 208.880 1416.300 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1399.120 208.880 1402.660 210.000 ;
  LAYER metal4 ;
  RECT 1399.120 208.880 1402.660 210.000 ;
  LAYER metal3 ;
  RECT 1399.120 208.880 1402.660 210.000 ;
  LAYER metal2 ;
  RECT 1399.120 208.880 1402.660 210.000 ;
  LAYER metal1 ;
  RECT 1399.120 208.880 1402.660 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1386.100 208.880 1389.640 210.000 ;
  LAYER metal4 ;
  RECT 1386.100 208.880 1389.640 210.000 ;
  LAYER metal3 ;
  RECT 1386.100 208.880 1389.640 210.000 ;
  LAYER metal2 ;
  RECT 1386.100 208.880 1389.640 210.000 ;
  LAYER metal1 ;
  RECT 1386.100 208.880 1389.640 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1372.460 208.880 1376.000 210.000 ;
  LAYER metal4 ;
  RECT 1372.460 208.880 1376.000 210.000 ;
  LAYER metal3 ;
  RECT 1372.460 208.880 1376.000 210.000 ;
  LAYER metal2 ;
  RECT 1372.460 208.880 1376.000 210.000 ;
  LAYER metal1 ;
  RECT 1372.460 208.880 1376.000 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1358.820 208.880 1362.360 210.000 ;
  LAYER metal4 ;
  RECT 1358.820 208.880 1362.360 210.000 ;
  LAYER metal3 ;
  RECT 1358.820 208.880 1362.360 210.000 ;
  LAYER metal2 ;
  RECT 1358.820 208.880 1362.360 210.000 ;
  LAYER metal1 ;
  RECT 1358.820 208.880 1362.360 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1291.860 208.880 1295.400 210.000 ;
  LAYER metal4 ;
  RECT 1291.860 208.880 1295.400 210.000 ;
  LAYER metal3 ;
  RECT 1291.860 208.880 1295.400 210.000 ;
  LAYER metal2 ;
  RECT 1291.860 208.880 1295.400 210.000 ;
  LAYER metal1 ;
  RECT 1291.860 208.880 1295.400 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1278.220 208.880 1281.760 210.000 ;
  LAYER metal4 ;
  RECT 1278.220 208.880 1281.760 210.000 ;
  LAYER metal3 ;
  RECT 1278.220 208.880 1281.760 210.000 ;
  LAYER metal2 ;
  RECT 1278.220 208.880 1281.760 210.000 ;
  LAYER metal1 ;
  RECT 1278.220 208.880 1281.760 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1264.580 208.880 1268.120 210.000 ;
  LAYER metal4 ;
  RECT 1264.580 208.880 1268.120 210.000 ;
  LAYER metal3 ;
  RECT 1264.580 208.880 1268.120 210.000 ;
  LAYER metal2 ;
  RECT 1264.580 208.880 1268.120 210.000 ;
  LAYER metal1 ;
  RECT 1264.580 208.880 1268.120 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1251.560 208.880 1255.100 210.000 ;
  LAYER metal4 ;
  RECT 1251.560 208.880 1255.100 210.000 ;
  LAYER metal3 ;
  RECT 1251.560 208.880 1255.100 210.000 ;
  LAYER metal2 ;
  RECT 1251.560 208.880 1255.100 210.000 ;
  LAYER metal1 ;
  RECT 1251.560 208.880 1255.100 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1237.920 208.880 1241.460 210.000 ;
  LAYER metal4 ;
  RECT 1237.920 208.880 1241.460 210.000 ;
  LAYER metal3 ;
  RECT 1237.920 208.880 1241.460 210.000 ;
  LAYER metal2 ;
  RECT 1237.920 208.880 1241.460 210.000 ;
  LAYER metal1 ;
  RECT 1237.920 208.880 1241.460 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1224.280 208.880 1227.820 210.000 ;
  LAYER metal4 ;
  RECT 1224.280 208.880 1227.820 210.000 ;
  LAYER metal3 ;
  RECT 1224.280 208.880 1227.820 210.000 ;
  LAYER metal2 ;
  RECT 1224.280 208.880 1227.820 210.000 ;
  LAYER metal1 ;
  RECT 1224.280 208.880 1227.820 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1157.320 208.880 1160.860 210.000 ;
  LAYER metal4 ;
  RECT 1157.320 208.880 1160.860 210.000 ;
  LAYER metal3 ;
  RECT 1157.320 208.880 1160.860 210.000 ;
  LAYER metal2 ;
  RECT 1157.320 208.880 1160.860 210.000 ;
  LAYER metal1 ;
  RECT 1157.320 208.880 1160.860 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1143.680 208.880 1147.220 210.000 ;
  LAYER metal4 ;
  RECT 1143.680 208.880 1147.220 210.000 ;
  LAYER metal3 ;
  RECT 1143.680 208.880 1147.220 210.000 ;
  LAYER metal2 ;
  RECT 1143.680 208.880 1147.220 210.000 ;
  LAYER metal1 ;
  RECT 1143.680 208.880 1147.220 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1130.660 208.880 1134.200 210.000 ;
  LAYER metal4 ;
  RECT 1130.660 208.880 1134.200 210.000 ;
  LAYER metal3 ;
  RECT 1130.660 208.880 1134.200 210.000 ;
  LAYER metal2 ;
  RECT 1130.660 208.880 1134.200 210.000 ;
  LAYER metal1 ;
  RECT 1130.660 208.880 1134.200 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1117.020 208.880 1120.560 210.000 ;
  LAYER metal4 ;
  RECT 1117.020 208.880 1120.560 210.000 ;
  LAYER metal3 ;
  RECT 1117.020 208.880 1120.560 210.000 ;
  LAYER metal2 ;
  RECT 1117.020 208.880 1120.560 210.000 ;
  LAYER metal1 ;
  RECT 1117.020 208.880 1120.560 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1103.380 208.880 1106.920 210.000 ;
  LAYER metal4 ;
  RECT 1103.380 208.880 1106.920 210.000 ;
  LAYER metal3 ;
  RECT 1103.380 208.880 1106.920 210.000 ;
  LAYER metal2 ;
  RECT 1103.380 208.880 1106.920 210.000 ;
  LAYER metal1 ;
  RECT 1103.380 208.880 1106.920 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1090.360 208.880 1093.900 210.000 ;
  LAYER metal4 ;
  RECT 1090.360 208.880 1093.900 210.000 ;
  LAYER metal3 ;
  RECT 1090.360 208.880 1093.900 210.000 ;
  LAYER metal2 ;
  RECT 1090.360 208.880 1093.900 210.000 ;
  LAYER metal1 ;
  RECT 1090.360 208.880 1093.900 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1022.780 208.880 1026.320 210.000 ;
  LAYER metal4 ;
  RECT 1022.780 208.880 1026.320 210.000 ;
  LAYER metal3 ;
  RECT 1022.780 208.880 1026.320 210.000 ;
  LAYER metal2 ;
  RECT 1022.780 208.880 1026.320 210.000 ;
  LAYER metal1 ;
  RECT 1022.780 208.880 1026.320 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1009.760 208.880 1013.300 210.000 ;
  LAYER metal4 ;
  RECT 1009.760 208.880 1013.300 210.000 ;
  LAYER metal3 ;
  RECT 1009.760 208.880 1013.300 210.000 ;
  LAYER metal2 ;
  RECT 1009.760 208.880 1013.300 210.000 ;
  LAYER metal1 ;
  RECT 1009.760 208.880 1013.300 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 996.120 208.880 999.660 210.000 ;
  LAYER metal4 ;
  RECT 996.120 208.880 999.660 210.000 ;
  LAYER metal3 ;
  RECT 996.120 208.880 999.660 210.000 ;
  LAYER metal2 ;
  RECT 996.120 208.880 999.660 210.000 ;
  LAYER metal1 ;
  RECT 996.120 208.880 999.660 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 982.480 208.880 986.020 210.000 ;
  LAYER metal4 ;
  RECT 982.480 208.880 986.020 210.000 ;
  LAYER metal3 ;
  RECT 982.480 208.880 986.020 210.000 ;
  LAYER metal2 ;
  RECT 982.480 208.880 986.020 210.000 ;
  LAYER metal1 ;
  RECT 982.480 208.880 986.020 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 969.460 208.880 973.000 210.000 ;
  LAYER metal4 ;
  RECT 969.460 208.880 973.000 210.000 ;
  LAYER metal3 ;
  RECT 969.460 208.880 973.000 210.000 ;
  LAYER metal2 ;
  RECT 969.460 208.880 973.000 210.000 ;
  LAYER metal1 ;
  RECT 969.460 208.880 973.000 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 955.820 208.880 959.360 210.000 ;
  LAYER metal4 ;
  RECT 955.820 208.880 959.360 210.000 ;
  LAYER metal3 ;
  RECT 955.820 208.880 959.360 210.000 ;
  LAYER metal2 ;
  RECT 955.820 208.880 959.360 210.000 ;
  LAYER metal1 ;
  RECT 955.820 208.880 959.360 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 888.240 208.880 891.780 210.000 ;
  LAYER metal4 ;
  RECT 888.240 208.880 891.780 210.000 ;
  LAYER metal3 ;
  RECT 888.240 208.880 891.780 210.000 ;
  LAYER metal2 ;
  RECT 888.240 208.880 891.780 210.000 ;
  LAYER metal1 ;
  RECT 888.240 208.880 891.780 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 875.220 208.880 878.760 210.000 ;
  LAYER metal4 ;
  RECT 875.220 208.880 878.760 210.000 ;
  LAYER metal3 ;
  RECT 875.220 208.880 878.760 210.000 ;
  LAYER metal2 ;
  RECT 875.220 208.880 878.760 210.000 ;
  LAYER metal1 ;
  RECT 875.220 208.880 878.760 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 861.580 208.880 865.120 210.000 ;
  LAYER metal4 ;
  RECT 861.580 208.880 865.120 210.000 ;
  LAYER metal3 ;
  RECT 861.580 208.880 865.120 210.000 ;
  LAYER metal2 ;
  RECT 861.580 208.880 865.120 210.000 ;
  LAYER metal1 ;
  RECT 861.580 208.880 865.120 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 847.940 208.880 851.480 210.000 ;
  LAYER metal4 ;
  RECT 847.940 208.880 851.480 210.000 ;
  LAYER metal3 ;
  RECT 847.940 208.880 851.480 210.000 ;
  LAYER metal2 ;
  RECT 847.940 208.880 851.480 210.000 ;
  LAYER metal1 ;
  RECT 847.940 208.880 851.480 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 834.920 208.880 838.460 210.000 ;
  LAYER metal4 ;
  RECT 834.920 208.880 838.460 210.000 ;
  LAYER metal3 ;
  RECT 834.920 208.880 838.460 210.000 ;
  LAYER metal2 ;
  RECT 834.920 208.880 838.460 210.000 ;
  LAYER metal1 ;
  RECT 834.920 208.880 838.460 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 821.280 208.880 824.820 210.000 ;
  LAYER metal4 ;
  RECT 821.280 208.880 824.820 210.000 ;
  LAYER metal3 ;
  RECT 821.280 208.880 824.820 210.000 ;
  LAYER metal2 ;
  RECT 821.280 208.880 824.820 210.000 ;
  LAYER metal1 ;
  RECT 821.280 208.880 824.820 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 754.320 208.880 757.860 210.000 ;
  LAYER metal4 ;
  RECT 754.320 208.880 757.860 210.000 ;
  LAYER metal3 ;
  RECT 754.320 208.880 757.860 210.000 ;
  LAYER metal2 ;
  RECT 754.320 208.880 757.860 210.000 ;
  LAYER metal1 ;
  RECT 754.320 208.880 757.860 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 740.680 208.880 744.220 210.000 ;
  LAYER metal4 ;
  RECT 740.680 208.880 744.220 210.000 ;
  LAYER metal3 ;
  RECT 740.680 208.880 744.220 210.000 ;
  LAYER metal2 ;
  RECT 740.680 208.880 744.220 210.000 ;
  LAYER metal1 ;
  RECT 740.680 208.880 744.220 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 727.040 208.880 730.580 210.000 ;
  LAYER metal4 ;
  RECT 727.040 208.880 730.580 210.000 ;
  LAYER metal3 ;
  RECT 727.040 208.880 730.580 210.000 ;
  LAYER metal2 ;
  RECT 727.040 208.880 730.580 210.000 ;
  LAYER metal1 ;
  RECT 727.040 208.880 730.580 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 714.020 208.880 717.560 210.000 ;
  LAYER metal4 ;
  RECT 714.020 208.880 717.560 210.000 ;
  LAYER metal3 ;
  RECT 714.020 208.880 717.560 210.000 ;
  LAYER metal2 ;
  RECT 714.020 208.880 717.560 210.000 ;
  LAYER metal1 ;
  RECT 714.020 208.880 717.560 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 700.380 208.880 703.920 210.000 ;
  LAYER metal4 ;
  RECT 700.380 208.880 703.920 210.000 ;
  LAYER metal3 ;
  RECT 700.380 208.880 703.920 210.000 ;
  LAYER metal2 ;
  RECT 700.380 208.880 703.920 210.000 ;
  LAYER metal1 ;
  RECT 700.380 208.880 703.920 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 686.740 208.880 690.280 210.000 ;
  LAYER metal4 ;
  RECT 686.740 208.880 690.280 210.000 ;
  LAYER metal3 ;
  RECT 686.740 208.880 690.280 210.000 ;
  LAYER metal2 ;
  RECT 686.740 208.880 690.280 210.000 ;
  LAYER metal1 ;
  RECT 686.740 208.880 690.280 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 619.780 208.880 623.320 210.000 ;
  LAYER metal4 ;
  RECT 619.780 208.880 623.320 210.000 ;
  LAYER metal3 ;
  RECT 619.780 208.880 623.320 210.000 ;
  LAYER metal2 ;
  RECT 619.780 208.880 623.320 210.000 ;
  LAYER metal1 ;
  RECT 619.780 208.880 623.320 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 606.140 208.880 609.680 210.000 ;
  LAYER metal4 ;
  RECT 606.140 208.880 609.680 210.000 ;
  LAYER metal3 ;
  RECT 606.140 208.880 609.680 210.000 ;
  LAYER metal2 ;
  RECT 606.140 208.880 609.680 210.000 ;
  LAYER metal1 ;
  RECT 606.140 208.880 609.680 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 593.120 208.880 596.660 210.000 ;
  LAYER metal4 ;
  RECT 593.120 208.880 596.660 210.000 ;
  LAYER metal3 ;
  RECT 593.120 208.880 596.660 210.000 ;
  LAYER metal2 ;
  RECT 593.120 208.880 596.660 210.000 ;
  LAYER metal1 ;
  RECT 593.120 208.880 596.660 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 579.480 208.880 583.020 210.000 ;
  LAYER metal4 ;
  RECT 579.480 208.880 583.020 210.000 ;
  LAYER metal3 ;
  RECT 579.480 208.880 583.020 210.000 ;
  LAYER metal2 ;
  RECT 579.480 208.880 583.020 210.000 ;
  LAYER metal1 ;
  RECT 579.480 208.880 583.020 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 565.840 208.880 569.380 210.000 ;
  LAYER metal4 ;
  RECT 565.840 208.880 569.380 210.000 ;
  LAYER metal3 ;
  RECT 565.840 208.880 569.380 210.000 ;
  LAYER metal2 ;
  RECT 565.840 208.880 569.380 210.000 ;
  LAYER metal1 ;
  RECT 565.840 208.880 569.380 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 552.820 208.880 556.360 210.000 ;
  LAYER metal4 ;
  RECT 552.820 208.880 556.360 210.000 ;
  LAYER metal3 ;
  RECT 552.820 208.880 556.360 210.000 ;
  LAYER metal2 ;
  RECT 552.820 208.880 556.360 210.000 ;
  LAYER metal1 ;
  RECT 552.820 208.880 556.360 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 485.240 208.880 488.780 210.000 ;
  LAYER metal4 ;
  RECT 485.240 208.880 488.780 210.000 ;
  LAYER metal3 ;
  RECT 485.240 208.880 488.780 210.000 ;
  LAYER metal2 ;
  RECT 485.240 208.880 488.780 210.000 ;
  LAYER metal1 ;
  RECT 485.240 208.880 488.780 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 471.600 208.880 475.140 210.000 ;
  LAYER metal4 ;
  RECT 471.600 208.880 475.140 210.000 ;
  LAYER metal3 ;
  RECT 471.600 208.880 475.140 210.000 ;
  LAYER metal2 ;
  RECT 471.600 208.880 475.140 210.000 ;
  LAYER metal1 ;
  RECT 471.600 208.880 475.140 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 458.580 208.880 462.120 210.000 ;
  LAYER metal4 ;
  RECT 458.580 208.880 462.120 210.000 ;
  LAYER metal3 ;
  RECT 458.580 208.880 462.120 210.000 ;
  LAYER metal2 ;
  RECT 458.580 208.880 462.120 210.000 ;
  LAYER metal1 ;
  RECT 458.580 208.880 462.120 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 444.940 208.880 448.480 210.000 ;
  LAYER metal4 ;
  RECT 444.940 208.880 448.480 210.000 ;
  LAYER metal3 ;
  RECT 444.940 208.880 448.480 210.000 ;
  LAYER metal2 ;
  RECT 444.940 208.880 448.480 210.000 ;
  LAYER metal1 ;
  RECT 444.940 208.880 448.480 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 431.300 208.880 434.840 210.000 ;
  LAYER metal4 ;
  RECT 431.300 208.880 434.840 210.000 ;
  LAYER metal3 ;
  RECT 431.300 208.880 434.840 210.000 ;
  LAYER metal2 ;
  RECT 431.300 208.880 434.840 210.000 ;
  LAYER metal1 ;
  RECT 431.300 208.880 434.840 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 418.280 208.880 421.820 210.000 ;
  LAYER metal4 ;
  RECT 418.280 208.880 421.820 210.000 ;
  LAYER metal3 ;
  RECT 418.280 208.880 421.820 210.000 ;
  LAYER metal2 ;
  RECT 418.280 208.880 421.820 210.000 ;
  LAYER metal1 ;
  RECT 418.280 208.880 421.820 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 350.700 208.880 354.240 210.000 ;
  LAYER metal4 ;
  RECT 350.700 208.880 354.240 210.000 ;
  LAYER metal3 ;
  RECT 350.700 208.880 354.240 210.000 ;
  LAYER metal2 ;
  RECT 350.700 208.880 354.240 210.000 ;
  LAYER metal1 ;
  RECT 350.700 208.880 354.240 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 337.680 208.880 341.220 210.000 ;
  LAYER metal4 ;
  RECT 337.680 208.880 341.220 210.000 ;
  LAYER metal3 ;
  RECT 337.680 208.880 341.220 210.000 ;
  LAYER metal2 ;
  RECT 337.680 208.880 341.220 210.000 ;
  LAYER metal1 ;
  RECT 337.680 208.880 341.220 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 324.040 208.880 327.580 210.000 ;
  LAYER metal4 ;
  RECT 324.040 208.880 327.580 210.000 ;
  LAYER metal3 ;
  RECT 324.040 208.880 327.580 210.000 ;
  LAYER metal2 ;
  RECT 324.040 208.880 327.580 210.000 ;
  LAYER metal1 ;
  RECT 324.040 208.880 327.580 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 310.400 208.880 313.940 210.000 ;
  LAYER metal4 ;
  RECT 310.400 208.880 313.940 210.000 ;
  LAYER metal3 ;
  RECT 310.400 208.880 313.940 210.000 ;
  LAYER metal2 ;
  RECT 310.400 208.880 313.940 210.000 ;
  LAYER metal1 ;
  RECT 310.400 208.880 313.940 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 297.380 208.880 300.920 210.000 ;
  LAYER metal4 ;
  RECT 297.380 208.880 300.920 210.000 ;
  LAYER metal3 ;
  RECT 297.380 208.880 300.920 210.000 ;
  LAYER metal2 ;
  RECT 297.380 208.880 300.920 210.000 ;
  LAYER metal1 ;
  RECT 297.380 208.880 300.920 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 283.740 208.880 287.280 210.000 ;
  LAYER metal4 ;
  RECT 283.740 208.880 287.280 210.000 ;
  LAYER metal3 ;
  RECT 283.740 208.880 287.280 210.000 ;
  LAYER metal2 ;
  RECT 283.740 208.880 287.280 210.000 ;
  LAYER metal1 ;
  RECT 283.740 208.880 287.280 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 216.780 208.880 220.320 210.000 ;
  LAYER metal4 ;
  RECT 216.780 208.880 220.320 210.000 ;
  LAYER metal3 ;
  RECT 216.780 208.880 220.320 210.000 ;
  LAYER metal2 ;
  RECT 216.780 208.880 220.320 210.000 ;
  LAYER metal1 ;
  RECT 216.780 208.880 220.320 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 203.140 208.880 206.680 210.000 ;
  LAYER metal4 ;
  RECT 203.140 208.880 206.680 210.000 ;
  LAYER metal3 ;
  RECT 203.140 208.880 206.680 210.000 ;
  LAYER metal2 ;
  RECT 203.140 208.880 206.680 210.000 ;
  LAYER metal1 ;
  RECT 203.140 208.880 206.680 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 189.500 208.880 193.040 210.000 ;
  LAYER metal4 ;
  RECT 189.500 208.880 193.040 210.000 ;
  LAYER metal3 ;
  RECT 189.500 208.880 193.040 210.000 ;
  LAYER metal2 ;
  RECT 189.500 208.880 193.040 210.000 ;
  LAYER metal1 ;
  RECT 189.500 208.880 193.040 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 176.480 208.880 180.020 210.000 ;
  LAYER metal4 ;
  RECT 176.480 208.880 180.020 210.000 ;
  LAYER metal3 ;
  RECT 176.480 208.880 180.020 210.000 ;
  LAYER metal2 ;
  RECT 176.480 208.880 180.020 210.000 ;
  LAYER metal1 ;
  RECT 176.480 208.880 180.020 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 162.840 208.880 166.380 210.000 ;
  LAYER metal4 ;
  RECT 162.840 208.880 166.380 210.000 ;
  LAYER metal3 ;
  RECT 162.840 208.880 166.380 210.000 ;
  LAYER metal2 ;
  RECT 162.840 208.880 166.380 210.000 ;
  LAYER metal1 ;
  RECT 162.840 208.880 166.380 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 149.200 208.880 152.740 210.000 ;
  LAYER metal4 ;
  RECT 149.200 208.880 152.740 210.000 ;
  LAYER metal3 ;
  RECT 149.200 208.880 152.740 210.000 ;
  LAYER metal2 ;
  RECT 149.200 208.880 152.740 210.000 ;
  LAYER metal1 ;
  RECT 149.200 208.880 152.740 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 82.240 208.880 85.780 210.000 ;
  LAYER metal4 ;
  RECT 82.240 208.880 85.780 210.000 ;
  LAYER metal3 ;
  RECT 82.240 208.880 85.780 210.000 ;
  LAYER metal2 ;
  RECT 82.240 208.880 85.780 210.000 ;
  LAYER metal1 ;
  RECT 82.240 208.880 85.780 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 68.600 208.880 72.140 210.000 ;
  LAYER metal4 ;
  RECT 68.600 208.880 72.140 210.000 ;
  LAYER metal3 ;
  RECT 68.600 208.880 72.140 210.000 ;
  LAYER metal2 ;
  RECT 68.600 208.880 72.140 210.000 ;
  LAYER metal1 ;
  RECT 68.600 208.880 72.140 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 54.960 208.880 58.500 210.000 ;
  LAYER metal4 ;
  RECT 54.960 208.880 58.500 210.000 ;
  LAYER metal3 ;
  RECT 54.960 208.880 58.500 210.000 ;
  LAYER metal2 ;
  RECT 54.960 208.880 58.500 210.000 ;
  LAYER metal1 ;
  RECT 54.960 208.880 58.500 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 41.940 208.880 45.480 210.000 ;
  LAYER metal4 ;
  RECT 41.940 208.880 45.480 210.000 ;
  LAYER metal3 ;
  RECT 41.940 208.880 45.480 210.000 ;
  LAYER metal2 ;
  RECT 41.940 208.880 45.480 210.000 ;
  LAYER metal1 ;
  RECT 41.940 208.880 45.480 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 28.300 208.880 31.840 210.000 ;
  LAYER metal4 ;
  RECT 28.300 208.880 31.840 210.000 ;
  LAYER metal3 ;
  RECT 28.300 208.880 31.840 210.000 ;
  LAYER metal2 ;
  RECT 28.300 208.880 31.840 210.000 ;
  LAYER metal1 ;
  RECT 28.300 208.880 31.840 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 14.660 208.880 18.200 210.000 ;
  LAYER metal4 ;
  RECT 14.660 208.880 18.200 210.000 ;
  LAYER metal3 ;
  RECT 14.660 208.880 18.200 210.000 ;
  LAYER metal2 ;
  RECT 14.660 208.880 18.200 210.000 ;
  LAYER metal1 ;
  RECT 14.660 208.880 18.200 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3555.480 0.000 3559.020 1.120 ;
  LAYER metal4 ;
  RECT 3555.480 0.000 3559.020 1.120 ;
  LAYER metal3 ;
  RECT 3555.480 0.000 3559.020 1.120 ;
  LAYER metal2 ;
  RECT 3555.480 0.000 3559.020 1.120 ;
  LAYER metal1 ;
  RECT 3555.480 0.000 3559.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3541.840 0.000 3545.380 1.120 ;
  LAYER metal4 ;
  RECT 3541.840 0.000 3545.380 1.120 ;
  LAYER metal3 ;
  RECT 3541.840 0.000 3545.380 1.120 ;
  LAYER metal2 ;
  RECT 3541.840 0.000 3545.380 1.120 ;
  LAYER metal1 ;
  RECT 3541.840 0.000 3545.380 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3528.820 0.000 3532.360 1.120 ;
  LAYER metal4 ;
  RECT 3528.820 0.000 3532.360 1.120 ;
  LAYER metal3 ;
  RECT 3528.820 0.000 3532.360 1.120 ;
  LAYER metal2 ;
  RECT 3528.820 0.000 3532.360 1.120 ;
  LAYER metal1 ;
  RECT 3528.820 0.000 3532.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3461.240 0.000 3464.780 1.120 ;
  LAYER metal4 ;
  RECT 3461.240 0.000 3464.780 1.120 ;
  LAYER metal3 ;
  RECT 3461.240 0.000 3464.780 1.120 ;
  LAYER metal2 ;
  RECT 3461.240 0.000 3464.780 1.120 ;
  LAYER metal1 ;
  RECT 3461.240 0.000 3464.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3447.600 0.000 3451.140 1.120 ;
  LAYER metal4 ;
  RECT 3447.600 0.000 3451.140 1.120 ;
  LAYER metal3 ;
  RECT 3447.600 0.000 3451.140 1.120 ;
  LAYER metal2 ;
  RECT 3447.600 0.000 3451.140 1.120 ;
  LAYER metal1 ;
  RECT 3447.600 0.000 3451.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3434.580 0.000 3438.120 1.120 ;
  LAYER metal4 ;
  RECT 3434.580 0.000 3438.120 1.120 ;
  LAYER metal3 ;
  RECT 3434.580 0.000 3438.120 1.120 ;
  LAYER metal2 ;
  RECT 3434.580 0.000 3438.120 1.120 ;
  LAYER metal1 ;
  RECT 3434.580 0.000 3438.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3420.940 0.000 3424.480 1.120 ;
  LAYER metal4 ;
  RECT 3420.940 0.000 3424.480 1.120 ;
  LAYER metal3 ;
  RECT 3420.940 0.000 3424.480 1.120 ;
  LAYER metal2 ;
  RECT 3420.940 0.000 3424.480 1.120 ;
  LAYER metal1 ;
  RECT 3420.940 0.000 3424.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3407.300 0.000 3410.840 1.120 ;
  LAYER metal4 ;
  RECT 3407.300 0.000 3410.840 1.120 ;
  LAYER metal3 ;
  RECT 3407.300 0.000 3410.840 1.120 ;
  LAYER metal2 ;
  RECT 3407.300 0.000 3410.840 1.120 ;
  LAYER metal1 ;
  RECT 3407.300 0.000 3410.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3394.280 0.000 3397.820 1.120 ;
  LAYER metal4 ;
  RECT 3394.280 0.000 3397.820 1.120 ;
  LAYER metal3 ;
  RECT 3394.280 0.000 3397.820 1.120 ;
  LAYER metal2 ;
  RECT 3394.280 0.000 3397.820 1.120 ;
  LAYER metal1 ;
  RECT 3394.280 0.000 3397.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3326.700 0.000 3330.240 1.120 ;
  LAYER metal4 ;
  RECT 3326.700 0.000 3330.240 1.120 ;
  LAYER metal3 ;
  RECT 3326.700 0.000 3330.240 1.120 ;
  LAYER metal2 ;
  RECT 3326.700 0.000 3330.240 1.120 ;
  LAYER metal1 ;
  RECT 3326.700 0.000 3330.240 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3313.680 0.000 3317.220 1.120 ;
  LAYER metal4 ;
  RECT 3313.680 0.000 3317.220 1.120 ;
  LAYER metal3 ;
  RECT 3313.680 0.000 3317.220 1.120 ;
  LAYER metal2 ;
  RECT 3313.680 0.000 3317.220 1.120 ;
  LAYER metal1 ;
  RECT 3313.680 0.000 3317.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3300.040 0.000 3303.580 1.120 ;
  LAYER metal4 ;
  RECT 3300.040 0.000 3303.580 1.120 ;
  LAYER metal3 ;
  RECT 3300.040 0.000 3303.580 1.120 ;
  LAYER metal2 ;
  RECT 3300.040 0.000 3303.580 1.120 ;
  LAYER metal1 ;
  RECT 3300.040 0.000 3303.580 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3286.400 0.000 3289.940 1.120 ;
  LAYER metal4 ;
  RECT 3286.400 0.000 3289.940 1.120 ;
  LAYER metal3 ;
  RECT 3286.400 0.000 3289.940 1.120 ;
  LAYER metal2 ;
  RECT 3286.400 0.000 3289.940 1.120 ;
  LAYER metal1 ;
  RECT 3286.400 0.000 3289.940 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3273.380 0.000 3276.920 1.120 ;
  LAYER metal4 ;
  RECT 3273.380 0.000 3276.920 1.120 ;
  LAYER metal3 ;
  RECT 3273.380 0.000 3276.920 1.120 ;
  LAYER metal2 ;
  RECT 3273.380 0.000 3276.920 1.120 ;
  LAYER metal1 ;
  RECT 3273.380 0.000 3276.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3259.740 0.000 3263.280 1.120 ;
  LAYER metal4 ;
  RECT 3259.740 0.000 3263.280 1.120 ;
  LAYER metal3 ;
  RECT 3259.740 0.000 3263.280 1.120 ;
  LAYER metal2 ;
  RECT 3259.740 0.000 3263.280 1.120 ;
  LAYER metal1 ;
  RECT 3259.740 0.000 3263.280 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3192.780 0.000 3196.320 1.120 ;
  LAYER metal4 ;
  RECT 3192.780 0.000 3196.320 1.120 ;
  LAYER metal3 ;
  RECT 3192.780 0.000 3196.320 1.120 ;
  LAYER metal2 ;
  RECT 3192.780 0.000 3196.320 1.120 ;
  LAYER metal1 ;
  RECT 3192.780 0.000 3196.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3179.140 0.000 3182.680 1.120 ;
  LAYER metal4 ;
  RECT 3179.140 0.000 3182.680 1.120 ;
  LAYER metal3 ;
  RECT 3179.140 0.000 3182.680 1.120 ;
  LAYER metal2 ;
  RECT 3179.140 0.000 3182.680 1.120 ;
  LAYER metal1 ;
  RECT 3179.140 0.000 3182.680 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3165.500 0.000 3169.040 1.120 ;
  LAYER metal4 ;
  RECT 3165.500 0.000 3169.040 1.120 ;
  LAYER metal3 ;
  RECT 3165.500 0.000 3169.040 1.120 ;
  LAYER metal2 ;
  RECT 3165.500 0.000 3169.040 1.120 ;
  LAYER metal1 ;
  RECT 3165.500 0.000 3169.040 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3152.480 0.000 3156.020 1.120 ;
  LAYER metal4 ;
  RECT 3152.480 0.000 3156.020 1.120 ;
  LAYER metal3 ;
  RECT 3152.480 0.000 3156.020 1.120 ;
  LAYER metal2 ;
  RECT 3152.480 0.000 3156.020 1.120 ;
  LAYER metal1 ;
  RECT 3152.480 0.000 3156.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3138.840 0.000 3142.380 1.120 ;
  LAYER metal4 ;
  RECT 3138.840 0.000 3142.380 1.120 ;
  LAYER metal3 ;
  RECT 3138.840 0.000 3142.380 1.120 ;
  LAYER metal2 ;
  RECT 3138.840 0.000 3142.380 1.120 ;
  LAYER metal1 ;
  RECT 3138.840 0.000 3142.380 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3125.200 0.000 3128.740 1.120 ;
  LAYER metal4 ;
  RECT 3125.200 0.000 3128.740 1.120 ;
  LAYER metal3 ;
  RECT 3125.200 0.000 3128.740 1.120 ;
  LAYER metal2 ;
  RECT 3125.200 0.000 3128.740 1.120 ;
  LAYER metal1 ;
  RECT 3125.200 0.000 3128.740 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3058.240 0.000 3061.780 1.120 ;
  LAYER metal4 ;
  RECT 3058.240 0.000 3061.780 1.120 ;
  LAYER metal3 ;
  RECT 3058.240 0.000 3061.780 1.120 ;
  LAYER metal2 ;
  RECT 3058.240 0.000 3061.780 1.120 ;
  LAYER metal1 ;
  RECT 3058.240 0.000 3061.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3044.600 0.000 3048.140 1.120 ;
  LAYER metal4 ;
  RECT 3044.600 0.000 3048.140 1.120 ;
  LAYER metal3 ;
  RECT 3044.600 0.000 3048.140 1.120 ;
  LAYER metal2 ;
  RECT 3044.600 0.000 3048.140 1.120 ;
  LAYER metal1 ;
  RECT 3044.600 0.000 3048.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3030.960 0.000 3034.500 1.120 ;
  LAYER metal4 ;
  RECT 3030.960 0.000 3034.500 1.120 ;
  LAYER metal3 ;
  RECT 3030.960 0.000 3034.500 1.120 ;
  LAYER metal2 ;
  RECT 3030.960 0.000 3034.500 1.120 ;
  LAYER metal1 ;
  RECT 3030.960 0.000 3034.500 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3017.940 0.000 3021.480 1.120 ;
  LAYER metal4 ;
  RECT 3017.940 0.000 3021.480 1.120 ;
  LAYER metal3 ;
  RECT 3017.940 0.000 3021.480 1.120 ;
  LAYER metal2 ;
  RECT 3017.940 0.000 3021.480 1.120 ;
  LAYER metal1 ;
  RECT 3017.940 0.000 3021.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3004.300 0.000 3007.840 1.120 ;
  LAYER metal4 ;
  RECT 3004.300 0.000 3007.840 1.120 ;
  LAYER metal3 ;
  RECT 3004.300 0.000 3007.840 1.120 ;
  LAYER metal2 ;
  RECT 3004.300 0.000 3007.840 1.120 ;
  LAYER metal1 ;
  RECT 3004.300 0.000 3007.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2990.660 0.000 2994.200 1.120 ;
  LAYER metal4 ;
  RECT 2990.660 0.000 2994.200 1.120 ;
  LAYER metal3 ;
  RECT 2990.660 0.000 2994.200 1.120 ;
  LAYER metal2 ;
  RECT 2990.660 0.000 2994.200 1.120 ;
  LAYER metal1 ;
  RECT 2990.660 0.000 2994.200 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2923.700 0.000 2927.240 1.120 ;
  LAYER metal4 ;
  RECT 2923.700 0.000 2927.240 1.120 ;
  LAYER metal3 ;
  RECT 2923.700 0.000 2927.240 1.120 ;
  LAYER metal2 ;
  RECT 2923.700 0.000 2927.240 1.120 ;
  LAYER metal1 ;
  RECT 2923.700 0.000 2927.240 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2910.060 0.000 2913.600 1.120 ;
  LAYER metal4 ;
  RECT 2910.060 0.000 2913.600 1.120 ;
  LAYER metal3 ;
  RECT 2910.060 0.000 2913.600 1.120 ;
  LAYER metal2 ;
  RECT 2910.060 0.000 2913.600 1.120 ;
  LAYER metal1 ;
  RECT 2910.060 0.000 2913.600 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2897.040 0.000 2900.580 1.120 ;
  LAYER metal4 ;
  RECT 2897.040 0.000 2900.580 1.120 ;
  LAYER metal3 ;
  RECT 2897.040 0.000 2900.580 1.120 ;
  LAYER metal2 ;
  RECT 2897.040 0.000 2900.580 1.120 ;
  LAYER metal1 ;
  RECT 2897.040 0.000 2900.580 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2883.400 0.000 2886.940 1.120 ;
  LAYER metal4 ;
  RECT 2883.400 0.000 2886.940 1.120 ;
  LAYER metal3 ;
  RECT 2883.400 0.000 2886.940 1.120 ;
  LAYER metal2 ;
  RECT 2883.400 0.000 2886.940 1.120 ;
  LAYER metal1 ;
  RECT 2883.400 0.000 2886.940 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2869.760 0.000 2873.300 1.120 ;
  LAYER metal4 ;
  RECT 2869.760 0.000 2873.300 1.120 ;
  LAYER metal3 ;
  RECT 2869.760 0.000 2873.300 1.120 ;
  LAYER metal2 ;
  RECT 2869.760 0.000 2873.300 1.120 ;
  LAYER metal1 ;
  RECT 2869.760 0.000 2873.300 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2856.740 0.000 2860.280 1.120 ;
  LAYER metal4 ;
  RECT 2856.740 0.000 2860.280 1.120 ;
  LAYER metal3 ;
  RECT 2856.740 0.000 2860.280 1.120 ;
  LAYER metal2 ;
  RECT 2856.740 0.000 2860.280 1.120 ;
  LAYER metal1 ;
  RECT 2856.740 0.000 2860.280 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2789.160 0.000 2792.700 1.120 ;
  LAYER metal4 ;
  RECT 2789.160 0.000 2792.700 1.120 ;
  LAYER metal3 ;
  RECT 2789.160 0.000 2792.700 1.120 ;
  LAYER metal2 ;
  RECT 2789.160 0.000 2792.700 1.120 ;
  LAYER metal1 ;
  RECT 2789.160 0.000 2792.700 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2776.140 0.000 2779.680 1.120 ;
  LAYER metal4 ;
  RECT 2776.140 0.000 2779.680 1.120 ;
  LAYER metal3 ;
  RECT 2776.140 0.000 2779.680 1.120 ;
  LAYER metal2 ;
  RECT 2776.140 0.000 2779.680 1.120 ;
  LAYER metal1 ;
  RECT 2776.140 0.000 2779.680 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2762.500 0.000 2766.040 1.120 ;
  LAYER metal4 ;
  RECT 2762.500 0.000 2766.040 1.120 ;
  LAYER metal3 ;
  RECT 2762.500 0.000 2766.040 1.120 ;
  LAYER metal2 ;
  RECT 2762.500 0.000 2766.040 1.120 ;
  LAYER metal1 ;
  RECT 2762.500 0.000 2766.040 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2748.860 0.000 2752.400 1.120 ;
  LAYER metal4 ;
  RECT 2748.860 0.000 2752.400 1.120 ;
  LAYER metal3 ;
  RECT 2748.860 0.000 2752.400 1.120 ;
  LAYER metal2 ;
  RECT 2748.860 0.000 2752.400 1.120 ;
  LAYER metal1 ;
  RECT 2748.860 0.000 2752.400 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2735.840 0.000 2739.380 1.120 ;
  LAYER metal4 ;
  RECT 2735.840 0.000 2739.380 1.120 ;
  LAYER metal3 ;
  RECT 2735.840 0.000 2739.380 1.120 ;
  LAYER metal2 ;
  RECT 2735.840 0.000 2739.380 1.120 ;
  LAYER metal1 ;
  RECT 2735.840 0.000 2739.380 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2722.200 0.000 2725.740 1.120 ;
  LAYER metal4 ;
  RECT 2722.200 0.000 2725.740 1.120 ;
  LAYER metal3 ;
  RECT 2722.200 0.000 2725.740 1.120 ;
  LAYER metal2 ;
  RECT 2722.200 0.000 2725.740 1.120 ;
  LAYER metal1 ;
  RECT 2722.200 0.000 2725.740 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2655.240 0.000 2658.780 1.120 ;
  LAYER metal4 ;
  RECT 2655.240 0.000 2658.780 1.120 ;
  LAYER metal3 ;
  RECT 2655.240 0.000 2658.780 1.120 ;
  LAYER metal2 ;
  RECT 2655.240 0.000 2658.780 1.120 ;
  LAYER metal1 ;
  RECT 2655.240 0.000 2658.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2641.600 0.000 2645.140 1.120 ;
  LAYER metal4 ;
  RECT 2641.600 0.000 2645.140 1.120 ;
  LAYER metal3 ;
  RECT 2641.600 0.000 2645.140 1.120 ;
  LAYER metal2 ;
  RECT 2641.600 0.000 2645.140 1.120 ;
  LAYER metal1 ;
  RECT 2641.600 0.000 2645.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2627.960 0.000 2631.500 1.120 ;
  LAYER metal4 ;
  RECT 2627.960 0.000 2631.500 1.120 ;
  LAYER metal3 ;
  RECT 2627.960 0.000 2631.500 1.120 ;
  LAYER metal2 ;
  RECT 2627.960 0.000 2631.500 1.120 ;
  LAYER metal1 ;
  RECT 2627.960 0.000 2631.500 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2614.320 0.000 2617.860 1.120 ;
  LAYER metal4 ;
  RECT 2614.320 0.000 2617.860 1.120 ;
  LAYER metal3 ;
  RECT 2614.320 0.000 2617.860 1.120 ;
  LAYER metal2 ;
  RECT 2614.320 0.000 2617.860 1.120 ;
  LAYER metal1 ;
  RECT 2614.320 0.000 2617.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2601.300 0.000 2604.840 1.120 ;
  LAYER metal4 ;
  RECT 2601.300 0.000 2604.840 1.120 ;
  LAYER metal3 ;
  RECT 2601.300 0.000 2604.840 1.120 ;
  LAYER metal2 ;
  RECT 2601.300 0.000 2604.840 1.120 ;
  LAYER metal1 ;
  RECT 2601.300 0.000 2604.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2587.660 0.000 2591.200 1.120 ;
  LAYER metal4 ;
  RECT 2587.660 0.000 2591.200 1.120 ;
  LAYER metal3 ;
  RECT 2587.660 0.000 2591.200 1.120 ;
  LAYER metal2 ;
  RECT 2587.660 0.000 2591.200 1.120 ;
  LAYER metal1 ;
  RECT 2587.660 0.000 2591.200 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2520.700 0.000 2524.240 1.120 ;
  LAYER metal4 ;
  RECT 2520.700 0.000 2524.240 1.120 ;
  LAYER metal3 ;
  RECT 2520.700 0.000 2524.240 1.120 ;
  LAYER metal2 ;
  RECT 2520.700 0.000 2524.240 1.120 ;
  LAYER metal1 ;
  RECT 2520.700 0.000 2524.240 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2507.060 0.000 2510.600 1.120 ;
  LAYER metal4 ;
  RECT 2507.060 0.000 2510.600 1.120 ;
  LAYER metal3 ;
  RECT 2507.060 0.000 2510.600 1.120 ;
  LAYER metal2 ;
  RECT 2507.060 0.000 2510.600 1.120 ;
  LAYER metal1 ;
  RECT 2507.060 0.000 2510.600 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2493.420 0.000 2496.960 1.120 ;
  LAYER metal4 ;
  RECT 2493.420 0.000 2496.960 1.120 ;
  LAYER metal3 ;
  RECT 2493.420 0.000 2496.960 1.120 ;
  LAYER metal2 ;
  RECT 2493.420 0.000 2496.960 1.120 ;
  LAYER metal1 ;
  RECT 2493.420 0.000 2496.960 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2480.400 0.000 2483.940 1.120 ;
  LAYER metal4 ;
  RECT 2480.400 0.000 2483.940 1.120 ;
  LAYER metal3 ;
  RECT 2480.400 0.000 2483.940 1.120 ;
  LAYER metal2 ;
  RECT 2480.400 0.000 2483.940 1.120 ;
  LAYER metal1 ;
  RECT 2480.400 0.000 2483.940 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2466.760 0.000 2470.300 1.120 ;
  LAYER metal4 ;
  RECT 2466.760 0.000 2470.300 1.120 ;
  LAYER metal3 ;
  RECT 2466.760 0.000 2470.300 1.120 ;
  LAYER metal2 ;
  RECT 2466.760 0.000 2470.300 1.120 ;
  LAYER metal1 ;
  RECT 2466.760 0.000 2470.300 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2453.120 0.000 2456.660 1.120 ;
  LAYER metal4 ;
  RECT 2453.120 0.000 2456.660 1.120 ;
  LAYER metal3 ;
  RECT 2453.120 0.000 2456.660 1.120 ;
  LAYER metal2 ;
  RECT 2453.120 0.000 2456.660 1.120 ;
  LAYER metal1 ;
  RECT 2453.120 0.000 2456.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2386.160 0.000 2389.700 1.120 ;
  LAYER metal4 ;
  RECT 2386.160 0.000 2389.700 1.120 ;
  LAYER metal3 ;
  RECT 2386.160 0.000 2389.700 1.120 ;
  LAYER metal2 ;
  RECT 2386.160 0.000 2389.700 1.120 ;
  LAYER metal1 ;
  RECT 2386.160 0.000 2389.700 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2372.520 0.000 2376.060 1.120 ;
  LAYER metal4 ;
  RECT 2372.520 0.000 2376.060 1.120 ;
  LAYER metal3 ;
  RECT 2372.520 0.000 2376.060 1.120 ;
  LAYER metal2 ;
  RECT 2372.520 0.000 2376.060 1.120 ;
  LAYER metal1 ;
  RECT 2372.520 0.000 2376.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2359.500 0.000 2363.040 1.120 ;
  LAYER metal4 ;
  RECT 2359.500 0.000 2363.040 1.120 ;
  LAYER metal3 ;
  RECT 2359.500 0.000 2363.040 1.120 ;
  LAYER metal2 ;
  RECT 2359.500 0.000 2363.040 1.120 ;
  LAYER metal1 ;
  RECT 2359.500 0.000 2363.040 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2345.860 0.000 2349.400 1.120 ;
  LAYER metal4 ;
  RECT 2345.860 0.000 2349.400 1.120 ;
  LAYER metal3 ;
  RECT 2345.860 0.000 2349.400 1.120 ;
  LAYER metal2 ;
  RECT 2345.860 0.000 2349.400 1.120 ;
  LAYER metal1 ;
  RECT 2345.860 0.000 2349.400 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2332.220 0.000 2335.760 1.120 ;
  LAYER metal4 ;
  RECT 2332.220 0.000 2335.760 1.120 ;
  LAYER metal3 ;
  RECT 2332.220 0.000 2335.760 1.120 ;
  LAYER metal2 ;
  RECT 2332.220 0.000 2335.760 1.120 ;
  LAYER metal1 ;
  RECT 2332.220 0.000 2335.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2319.200 0.000 2322.740 1.120 ;
  LAYER metal4 ;
  RECT 2319.200 0.000 2322.740 1.120 ;
  LAYER metal3 ;
  RECT 2319.200 0.000 2322.740 1.120 ;
  LAYER metal2 ;
  RECT 2319.200 0.000 2322.740 1.120 ;
  LAYER metal1 ;
  RECT 2319.200 0.000 2322.740 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2251.620 0.000 2255.160 1.120 ;
  LAYER metal4 ;
  RECT 2251.620 0.000 2255.160 1.120 ;
  LAYER metal3 ;
  RECT 2251.620 0.000 2255.160 1.120 ;
  LAYER metal2 ;
  RECT 2251.620 0.000 2255.160 1.120 ;
  LAYER metal1 ;
  RECT 2251.620 0.000 2255.160 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2238.600 0.000 2242.140 1.120 ;
  LAYER metal4 ;
  RECT 2238.600 0.000 2242.140 1.120 ;
  LAYER metal3 ;
  RECT 2238.600 0.000 2242.140 1.120 ;
  LAYER metal2 ;
  RECT 2238.600 0.000 2242.140 1.120 ;
  LAYER metal1 ;
  RECT 2238.600 0.000 2242.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2224.960 0.000 2228.500 1.120 ;
  LAYER metal4 ;
  RECT 2224.960 0.000 2228.500 1.120 ;
  LAYER metal3 ;
  RECT 2224.960 0.000 2228.500 1.120 ;
  LAYER metal2 ;
  RECT 2224.960 0.000 2228.500 1.120 ;
  LAYER metal1 ;
  RECT 2224.960 0.000 2228.500 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2211.320 0.000 2214.860 1.120 ;
  LAYER metal4 ;
  RECT 2211.320 0.000 2214.860 1.120 ;
  LAYER metal3 ;
  RECT 2211.320 0.000 2214.860 1.120 ;
  LAYER metal2 ;
  RECT 2211.320 0.000 2214.860 1.120 ;
  LAYER metal1 ;
  RECT 2211.320 0.000 2214.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2197.680 0.000 2201.220 1.120 ;
  LAYER metal4 ;
  RECT 2197.680 0.000 2201.220 1.120 ;
  LAYER metal3 ;
  RECT 2197.680 0.000 2201.220 1.120 ;
  LAYER metal2 ;
  RECT 2197.680 0.000 2201.220 1.120 ;
  LAYER metal1 ;
  RECT 2197.680 0.000 2201.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2184.660 0.000 2188.200 1.120 ;
  LAYER metal4 ;
  RECT 2184.660 0.000 2188.200 1.120 ;
  LAYER metal3 ;
  RECT 2184.660 0.000 2188.200 1.120 ;
  LAYER metal2 ;
  RECT 2184.660 0.000 2188.200 1.120 ;
  LAYER metal1 ;
  RECT 2184.660 0.000 2188.200 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2117.080 0.000 2120.620 1.120 ;
  LAYER metal4 ;
  RECT 2117.080 0.000 2120.620 1.120 ;
  LAYER metal3 ;
  RECT 2117.080 0.000 2120.620 1.120 ;
  LAYER metal2 ;
  RECT 2117.080 0.000 2120.620 1.120 ;
  LAYER metal1 ;
  RECT 2117.080 0.000 2120.620 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2104.060 0.000 2107.600 1.120 ;
  LAYER metal4 ;
  RECT 2104.060 0.000 2107.600 1.120 ;
  LAYER metal3 ;
  RECT 2104.060 0.000 2107.600 1.120 ;
  LAYER metal2 ;
  RECT 2104.060 0.000 2107.600 1.120 ;
  LAYER metal1 ;
  RECT 2104.060 0.000 2107.600 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2090.420 0.000 2093.960 1.120 ;
  LAYER metal4 ;
  RECT 2090.420 0.000 2093.960 1.120 ;
  LAYER metal3 ;
  RECT 2090.420 0.000 2093.960 1.120 ;
  LAYER metal2 ;
  RECT 2090.420 0.000 2093.960 1.120 ;
  LAYER metal1 ;
  RECT 2090.420 0.000 2093.960 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2076.780 0.000 2080.320 1.120 ;
  LAYER metal4 ;
  RECT 2076.780 0.000 2080.320 1.120 ;
  LAYER metal3 ;
  RECT 2076.780 0.000 2080.320 1.120 ;
  LAYER metal2 ;
  RECT 2076.780 0.000 2080.320 1.120 ;
  LAYER metal1 ;
  RECT 2076.780 0.000 2080.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2063.760 0.000 2067.300 1.120 ;
  LAYER metal4 ;
  RECT 2063.760 0.000 2067.300 1.120 ;
  LAYER metal3 ;
  RECT 2063.760 0.000 2067.300 1.120 ;
  LAYER metal2 ;
  RECT 2063.760 0.000 2067.300 1.120 ;
  LAYER metal1 ;
  RECT 2063.760 0.000 2067.300 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2050.120 0.000 2053.660 1.120 ;
  LAYER metal4 ;
  RECT 2050.120 0.000 2053.660 1.120 ;
  LAYER metal3 ;
  RECT 2050.120 0.000 2053.660 1.120 ;
  LAYER metal2 ;
  RECT 2050.120 0.000 2053.660 1.120 ;
  LAYER metal1 ;
  RECT 2050.120 0.000 2053.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1983.160 0.000 1986.700 1.120 ;
  LAYER metal4 ;
  RECT 1983.160 0.000 1986.700 1.120 ;
  LAYER metal3 ;
  RECT 1983.160 0.000 1986.700 1.120 ;
  LAYER metal2 ;
  RECT 1983.160 0.000 1986.700 1.120 ;
  LAYER metal1 ;
  RECT 1983.160 0.000 1986.700 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1969.520 0.000 1973.060 1.120 ;
  LAYER metal4 ;
  RECT 1969.520 0.000 1973.060 1.120 ;
  LAYER metal3 ;
  RECT 1969.520 0.000 1973.060 1.120 ;
  LAYER metal2 ;
  RECT 1969.520 0.000 1973.060 1.120 ;
  LAYER metal1 ;
  RECT 1969.520 0.000 1973.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1955.880 0.000 1959.420 1.120 ;
  LAYER metal4 ;
  RECT 1955.880 0.000 1959.420 1.120 ;
  LAYER metal3 ;
  RECT 1955.880 0.000 1959.420 1.120 ;
  LAYER metal2 ;
  RECT 1955.880 0.000 1959.420 1.120 ;
  LAYER metal1 ;
  RECT 1955.880 0.000 1959.420 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1942.860 0.000 1946.400 1.120 ;
  LAYER metal4 ;
  RECT 1942.860 0.000 1946.400 1.120 ;
  LAYER metal3 ;
  RECT 1942.860 0.000 1946.400 1.120 ;
  LAYER metal2 ;
  RECT 1942.860 0.000 1946.400 1.120 ;
  LAYER metal1 ;
  RECT 1942.860 0.000 1946.400 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1929.220 0.000 1932.760 1.120 ;
  LAYER metal4 ;
  RECT 1929.220 0.000 1932.760 1.120 ;
  LAYER metal3 ;
  RECT 1929.220 0.000 1932.760 1.120 ;
  LAYER metal2 ;
  RECT 1929.220 0.000 1932.760 1.120 ;
  LAYER metal1 ;
  RECT 1929.220 0.000 1932.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1915.580 0.000 1919.120 1.120 ;
  LAYER metal4 ;
  RECT 1915.580 0.000 1919.120 1.120 ;
  LAYER metal3 ;
  RECT 1915.580 0.000 1919.120 1.120 ;
  LAYER metal2 ;
  RECT 1915.580 0.000 1919.120 1.120 ;
  LAYER metal1 ;
  RECT 1915.580 0.000 1919.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1848.620 0.000 1852.160 1.120 ;
  LAYER metal4 ;
  RECT 1848.620 0.000 1852.160 1.120 ;
  LAYER metal3 ;
  RECT 1848.620 0.000 1852.160 1.120 ;
  LAYER metal2 ;
  RECT 1848.620 0.000 1852.160 1.120 ;
  LAYER metal1 ;
  RECT 1848.620 0.000 1852.160 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1834.980 0.000 1838.520 1.120 ;
  LAYER metal4 ;
  RECT 1834.980 0.000 1838.520 1.120 ;
  LAYER metal3 ;
  RECT 1834.980 0.000 1838.520 1.120 ;
  LAYER metal2 ;
  RECT 1834.980 0.000 1838.520 1.120 ;
  LAYER metal1 ;
  RECT 1834.980 0.000 1838.520 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1826.300 0.000 1829.840 1.120 ;
  LAYER metal4 ;
  RECT 1826.300 0.000 1829.840 1.120 ;
  LAYER metal3 ;
  RECT 1826.300 0.000 1829.840 1.120 ;
  LAYER metal2 ;
  RECT 1826.300 0.000 1829.840 1.120 ;
  LAYER metal1 ;
  RECT 1826.300 0.000 1829.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1817.620 0.000 1821.160 1.120 ;
  LAYER metal4 ;
  RECT 1817.620 0.000 1821.160 1.120 ;
  LAYER metal3 ;
  RECT 1817.620 0.000 1821.160 1.120 ;
  LAYER metal2 ;
  RECT 1817.620 0.000 1821.160 1.120 ;
  LAYER metal1 ;
  RECT 1817.620 0.000 1821.160 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1803.980 0.000 1807.520 1.120 ;
  LAYER metal4 ;
  RECT 1803.980 0.000 1807.520 1.120 ;
  LAYER metal3 ;
  RECT 1803.980 0.000 1807.520 1.120 ;
  LAYER metal2 ;
  RECT 1803.980 0.000 1807.520 1.120 ;
  LAYER metal1 ;
  RECT 1803.980 0.000 1807.520 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1758.720 0.000 1762.260 1.120 ;
  LAYER metal4 ;
  RECT 1758.720 0.000 1762.260 1.120 ;
  LAYER metal3 ;
  RECT 1758.720 0.000 1762.260 1.120 ;
  LAYER metal2 ;
  RECT 1758.720 0.000 1762.260 1.120 ;
  LAYER metal1 ;
  RECT 1758.720 0.000 1762.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1694.860 0.000 1698.400 1.120 ;
  LAYER metal4 ;
  RECT 1694.860 0.000 1698.400 1.120 ;
  LAYER metal3 ;
  RECT 1694.860 0.000 1698.400 1.120 ;
  LAYER metal2 ;
  RECT 1694.860 0.000 1698.400 1.120 ;
  LAYER metal1 ;
  RECT 1694.860 0.000 1698.400 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1681.220 0.000 1684.760 1.120 ;
  LAYER metal4 ;
  RECT 1681.220 0.000 1684.760 1.120 ;
  LAYER metal3 ;
  RECT 1681.220 0.000 1684.760 1.120 ;
  LAYER metal2 ;
  RECT 1681.220 0.000 1684.760 1.120 ;
  LAYER metal1 ;
  RECT 1681.220 0.000 1684.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1668.200 0.000 1671.740 1.120 ;
  LAYER metal4 ;
  RECT 1668.200 0.000 1671.740 1.120 ;
  LAYER metal3 ;
  RECT 1668.200 0.000 1671.740 1.120 ;
  LAYER metal2 ;
  RECT 1668.200 0.000 1671.740 1.120 ;
  LAYER metal1 ;
  RECT 1668.200 0.000 1671.740 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1654.560 0.000 1658.100 1.120 ;
  LAYER metal4 ;
  RECT 1654.560 0.000 1658.100 1.120 ;
  LAYER metal3 ;
  RECT 1654.560 0.000 1658.100 1.120 ;
  LAYER metal2 ;
  RECT 1654.560 0.000 1658.100 1.120 ;
  LAYER metal1 ;
  RECT 1654.560 0.000 1658.100 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1640.920 0.000 1644.460 1.120 ;
  LAYER metal4 ;
  RECT 1640.920 0.000 1644.460 1.120 ;
  LAYER metal3 ;
  RECT 1640.920 0.000 1644.460 1.120 ;
  LAYER metal2 ;
  RECT 1640.920 0.000 1644.460 1.120 ;
  LAYER metal1 ;
  RECT 1640.920 0.000 1644.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1627.900 0.000 1631.440 1.120 ;
  LAYER metal4 ;
  RECT 1627.900 0.000 1631.440 1.120 ;
  LAYER metal3 ;
  RECT 1627.900 0.000 1631.440 1.120 ;
  LAYER metal2 ;
  RECT 1627.900 0.000 1631.440 1.120 ;
  LAYER metal1 ;
  RECT 1627.900 0.000 1631.440 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1560.320 0.000 1563.860 1.120 ;
  LAYER metal4 ;
  RECT 1560.320 0.000 1563.860 1.120 ;
  LAYER metal3 ;
  RECT 1560.320 0.000 1563.860 1.120 ;
  LAYER metal2 ;
  RECT 1560.320 0.000 1563.860 1.120 ;
  LAYER metal1 ;
  RECT 1560.320 0.000 1563.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1547.300 0.000 1550.840 1.120 ;
  LAYER metal4 ;
  RECT 1547.300 0.000 1550.840 1.120 ;
  LAYER metal3 ;
  RECT 1547.300 0.000 1550.840 1.120 ;
  LAYER metal2 ;
  RECT 1547.300 0.000 1550.840 1.120 ;
  LAYER metal1 ;
  RECT 1547.300 0.000 1550.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1533.660 0.000 1537.200 1.120 ;
  LAYER metal4 ;
  RECT 1533.660 0.000 1537.200 1.120 ;
  LAYER metal3 ;
  RECT 1533.660 0.000 1537.200 1.120 ;
  LAYER metal2 ;
  RECT 1533.660 0.000 1537.200 1.120 ;
  LAYER metal1 ;
  RECT 1533.660 0.000 1537.200 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1520.020 0.000 1523.560 1.120 ;
  LAYER metal4 ;
  RECT 1520.020 0.000 1523.560 1.120 ;
  LAYER metal3 ;
  RECT 1520.020 0.000 1523.560 1.120 ;
  LAYER metal2 ;
  RECT 1520.020 0.000 1523.560 1.120 ;
  LAYER metal1 ;
  RECT 1520.020 0.000 1523.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1507.000 0.000 1510.540 1.120 ;
  LAYER metal4 ;
  RECT 1507.000 0.000 1510.540 1.120 ;
  LAYER metal3 ;
  RECT 1507.000 0.000 1510.540 1.120 ;
  LAYER metal2 ;
  RECT 1507.000 0.000 1510.540 1.120 ;
  LAYER metal1 ;
  RECT 1507.000 0.000 1510.540 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1493.360 0.000 1496.900 1.120 ;
  LAYER metal4 ;
  RECT 1493.360 0.000 1496.900 1.120 ;
  LAYER metal3 ;
  RECT 1493.360 0.000 1496.900 1.120 ;
  LAYER metal2 ;
  RECT 1493.360 0.000 1496.900 1.120 ;
  LAYER metal1 ;
  RECT 1493.360 0.000 1496.900 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1426.400 0.000 1429.940 1.120 ;
  LAYER metal4 ;
  RECT 1426.400 0.000 1429.940 1.120 ;
  LAYER metal3 ;
  RECT 1426.400 0.000 1429.940 1.120 ;
  LAYER metal2 ;
  RECT 1426.400 0.000 1429.940 1.120 ;
  LAYER metal1 ;
  RECT 1426.400 0.000 1429.940 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1412.760 0.000 1416.300 1.120 ;
  LAYER metal4 ;
  RECT 1412.760 0.000 1416.300 1.120 ;
  LAYER metal3 ;
  RECT 1412.760 0.000 1416.300 1.120 ;
  LAYER metal2 ;
  RECT 1412.760 0.000 1416.300 1.120 ;
  LAYER metal1 ;
  RECT 1412.760 0.000 1416.300 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1399.120 0.000 1402.660 1.120 ;
  LAYER metal4 ;
  RECT 1399.120 0.000 1402.660 1.120 ;
  LAYER metal3 ;
  RECT 1399.120 0.000 1402.660 1.120 ;
  LAYER metal2 ;
  RECT 1399.120 0.000 1402.660 1.120 ;
  LAYER metal1 ;
  RECT 1399.120 0.000 1402.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1386.100 0.000 1389.640 1.120 ;
  LAYER metal4 ;
  RECT 1386.100 0.000 1389.640 1.120 ;
  LAYER metal3 ;
  RECT 1386.100 0.000 1389.640 1.120 ;
  LAYER metal2 ;
  RECT 1386.100 0.000 1389.640 1.120 ;
  LAYER metal1 ;
  RECT 1386.100 0.000 1389.640 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1372.460 0.000 1376.000 1.120 ;
  LAYER metal4 ;
  RECT 1372.460 0.000 1376.000 1.120 ;
  LAYER metal3 ;
  RECT 1372.460 0.000 1376.000 1.120 ;
  LAYER metal2 ;
  RECT 1372.460 0.000 1376.000 1.120 ;
  LAYER metal1 ;
  RECT 1372.460 0.000 1376.000 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1358.820 0.000 1362.360 1.120 ;
  LAYER metal4 ;
  RECT 1358.820 0.000 1362.360 1.120 ;
  LAYER metal3 ;
  RECT 1358.820 0.000 1362.360 1.120 ;
  LAYER metal2 ;
  RECT 1358.820 0.000 1362.360 1.120 ;
  LAYER metal1 ;
  RECT 1358.820 0.000 1362.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1291.860 0.000 1295.400 1.120 ;
  LAYER metal4 ;
  RECT 1291.860 0.000 1295.400 1.120 ;
  LAYER metal3 ;
  RECT 1291.860 0.000 1295.400 1.120 ;
  LAYER metal2 ;
  RECT 1291.860 0.000 1295.400 1.120 ;
  LAYER metal1 ;
  RECT 1291.860 0.000 1295.400 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1278.220 0.000 1281.760 1.120 ;
  LAYER metal4 ;
  RECT 1278.220 0.000 1281.760 1.120 ;
  LAYER metal3 ;
  RECT 1278.220 0.000 1281.760 1.120 ;
  LAYER metal2 ;
  RECT 1278.220 0.000 1281.760 1.120 ;
  LAYER metal1 ;
  RECT 1278.220 0.000 1281.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1264.580 0.000 1268.120 1.120 ;
  LAYER metal4 ;
  RECT 1264.580 0.000 1268.120 1.120 ;
  LAYER metal3 ;
  RECT 1264.580 0.000 1268.120 1.120 ;
  LAYER metal2 ;
  RECT 1264.580 0.000 1268.120 1.120 ;
  LAYER metal1 ;
  RECT 1264.580 0.000 1268.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1251.560 0.000 1255.100 1.120 ;
  LAYER metal4 ;
  RECT 1251.560 0.000 1255.100 1.120 ;
  LAYER metal3 ;
  RECT 1251.560 0.000 1255.100 1.120 ;
  LAYER metal2 ;
  RECT 1251.560 0.000 1255.100 1.120 ;
  LAYER metal1 ;
  RECT 1251.560 0.000 1255.100 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1237.920 0.000 1241.460 1.120 ;
  LAYER metal4 ;
  RECT 1237.920 0.000 1241.460 1.120 ;
  LAYER metal3 ;
  RECT 1237.920 0.000 1241.460 1.120 ;
  LAYER metal2 ;
  RECT 1237.920 0.000 1241.460 1.120 ;
  LAYER metal1 ;
  RECT 1237.920 0.000 1241.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1224.280 0.000 1227.820 1.120 ;
  LAYER metal4 ;
  RECT 1224.280 0.000 1227.820 1.120 ;
  LAYER metal3 ;
  RECT 1224.280 0.000 1227.820 1.120 ;
  LAYER metal2 ;
  RECT 1224.280 0.000 1227.820 1.120 ;
  LAYER metal1 ;
  RECT 1224.280 0.000 1227.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1157.320 0.000 1160.860 1.120 ;
  LAYER metal4 ;
  RECT 1157.320 0.000 1160.860 1.120 ;
  LAYER metal3 ;
  RECT 1157.320 0.000 1160.860 1.120 ;
  LAYER metal2 ;
  RECT 1157.320 0.000 1160.860 1.120 ;
  LAYER metal1 ;
  RECT 1157.320 0.000 1160.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1143.680 0.000 1147.220 1.120 ;
  LAYER metal4 ;
  RECT 1143.680 0.000 1147.220 1.120 ;
  LAYER metal3 ;
  RECT 1143.680 0.000 1147.220 1.120 ;
  LAYER metal2 ;
  RECT 1143.680 0.000 1147.220 1.120 ;
  LAYER metal1 ;
  RECT 1143.680 0.000 1147.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1130.660 0.000 1134.200 1.120 ;
  LAYER metal4 ;
  RECT 1130.660 0.000 1134.200 1.120 ;
  LAYER metal3 ;
  RECT 1130.660 0.000 1134.200 1.120 ;
  LAYER metal2 ;
  RECT 1130.660 0.000 1134.200 1.120 ;
  LAYER metal1 ;
  RECT 1130.660 0.000 1134.200 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1117.020 0.000 1120.560 1.120 ;
  LAYER metal4 ;
  RECT 1117.020 0.000 1120.560 1.120 ;
  LAYER metal3 ;
  RECT 1117.020 0.000 1120.560 1.120 ;
  LAYER metal2 ;
  RECT 1117.020 0.000 1120.560 1.120 ;
  LAYER metal1 ;
  RECT 1117.020 0.000 1120.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1103.380 0.000 1106.920 1.120 ;
  LAYER metal4 ;
  RECT 1103.380 0.000 1106.920 1.120 ;
  LAYER metal3 ;
  RECT 1103.380 0.000 1106.920 1.120 ;
  LAYER metal2 ;
  RECT 1103.380 0.000 1106.920 1.120 ;
  LAYER metal1 ;
  RECT 1103.380 0.000 1106.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1090.360 0.000 1093.900 1.120 ;
  LAYER metal4 ;
  RECT 1090.360 0.000 1093.900 1.120 ;
  LAYER metal3 ;
  RECT 1090.360 0.000 1093.900 1.120 ;
  LAYER metal2 ;
  RECT 1090.360 0.000 1093.900 1.120 ;
  LAYER metal1 ;
  RECT 1090.360 0.000 1093.900 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1022.780 0.000 1026.320 1.120 ;
  LAYER metal4 ;
  RECT 1022.780 0.000 1026.320 1.120 ;
  LAYER metal3 ;
  RECT 1022.780 0.000 1026.320 1.120 ;
  LAYER metal2 ;
  RECT 1022.780 0.000 1026.320 1.120 ;
  LAYER metal1 ;
  RECT 1022.780 0.000 1026.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1009.760 0.000 1013.300 1.120 ;
  LAYER metal4 ;
  RECT 1009.760 0.000 1013.300 1.120 ;
  LAYER metal3 ;
  RECT 1009.760 0.000 1013.300 1.120 ;
  LAYER metal2 ;
  RECT 1009.760 0.000 1013.300 1.120 ;
  LAYER metal1 ;
  RECT 1009.760 0.000 1013.300 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 996.120 0.000 999.660 1.120 ;
  LAYER metal4 ;
  RECT 996.120 0.000 999.660 1.120 ;
  LAYER metal3 ;
  RECT 996.120 0.000 999.660 1.120 ;
  LAYER metal2 ;
  RECT 996.120 0.000 999.660 1.120 ;
  LAYER metal1 ;
  RECT 996.120 0.000 999.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 982.480 0.000 986.020 1.120 ;
  LAYER metal4 ;
  RECT 982.480 0.000 986.020 1.120 ;
  LAYER metal3 ;
  RECT 982.480 0.000 986.020 1.120 ;
  LAYER metal2 ;
  RECT 982.480 0.000 986.020 1.120 ;
  LAYER metal1 ;
  RECT 982.480 0.000 986.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 969.460 0.000 973.000 1.120 ;
  LAYER metal4 ;
  RECT 969.460 0.000 973.000 1.120 ;
  LAYER metal3 ;
  RECT 969.460 0.000 973.000 1.120 ;
  LAYER metal2 ;
  RECT 969.460 0.000 973.000 1.120 ;
  LAYER metal1 ;
  RECT 969.460 0.000 973.000 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 955.820 0.000 959.360 1.120 ;
  LAYER metal4 ;
  RECT 955.820 0.000 959.360 1.120 ;
  LAYER metal3 ;
  RECT 955.820 0.000 959.360 1.120 ;
  LAYER metal2 ;
  RECT 955.820 0.000 959.360 1.120 ;
  LAYER metal1 ;
  RECT 955.820 0.000 959.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 888.240 0.000 891.780 1.120 ;
  LAYER metal4 ;
  RECT 888.240 0.000 891.780 1.120 ;
  LAYER metal3 ;
  RECT 888.240 0.000 891.780 1.120 ;
  LAYER metal2 ;
  RECT 888.240 0.000 891.780 1.120 ;
  LAYER metal1 ;
  RECT 888.240 0.000 891.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 875.220 0.000 878.760 1.120 ;
  LAYER metal4 ;
  RECT 875.220 0.000 878.760 1.120 ;
  LAYER metal3 ;
  RECT 875.220 0.000 878.760 1.120 ;
  LAYER metal2 ;
  RECT 875.220 0.000 878.760 1.120 ;
  LAYER metal1 ;
  RECT 875.220 0.000 878.760 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 861.580 0.000 865.120 1.120 ;
  LAYER metal4 ;
  RECT 861.580 0.000 865.120 1.120 ;
  LAYER metal3 ;
  RECT 861.580 0.000 865.120 1.120 ;
  LAYER metal2 ;
  RECT 861.580 0.000 865.120 1.120 ;
  LAYER metal1 ;
  RECT 861.580 0.000 865.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 847.940 0.000 851.480 1.120 ;
  LAYER metal4 ;
  RECT 847.940 0.000 851.480 1.120 ;
  LAYER metal3 ;
  RECT 847.940 0.000 851.480 1.120 ;
  LAYER metal2 ;
  RECT 847.940 0.000 851.480 1.120 ;
  LAYER metal1 ;
  RECT 847.940 0.000 851.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 834.920 0.000 838.460 1.120 ;
  LAYER metal4 ;
  RECT 834.920 0.000 838.460 1.120 ;
  LAYER metal3 ;
  RECT 834.920 0.000 838.460 1.120 ;
  LAYER metal2 ;
  RECT 834.920 0.000 838.460 1.120 ;
  LAYER metal1 ;
  RECT 834.920 0.000 838.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 821.280 0.000 824.820 1.120 ;
  LAYER metal4 ;
  RECT 821.280 0.000 824.820 1.120 ;
  LAYER metal3 ;
  RECT 821.280 0.000 824.820 1.120 ;
  LAYER metal2 ;
  RECT 821.280 0.000 824.820 1.120 ;
  LAYER metal1 ;
  RECT 821.280 0.000 824.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 754.320 0.000 757.860 1.120 ;
  LAYER metal4 ;
  RECT 754.320 0.000 757.860 1.120 ;
  LAYER metal3 ;
  RECT 754.320 0.000 757.860 1.120 ;
  LAYER metal2 ;
  RECT 754.320 0.000 757.860 1.120 ;
  LAYER metal1 ;
  RECT 754.320 0.000 757.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 740.680 0.000 744.220 1.120 ;
  LAYER metal4 ;
  RECT 740.680 0.000 744.220 1.120 ;
  LAYER metal3 ;
  RECT 740.680 0.000 744.220 1.120 ;
  LAYER metal2 ;
  RECT 740.680 0.000 744.220 1.120 ;
  LAYER metal1 ;
  RECT 740.680 0.000 744.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 727.040 0.000 730.580 1.120 ;
  LAYER metal4 ;
  RECT 727.040 0.000 730.580 1.120 ;
  LAYER metal3 ;
  RECT 727.040 0.000 730.580 1.120 ;
  LAYER metal2 ;
  RECT 727.040 0.000 730.580 1.120 ;
  LAYER metal1 ;
  RECT 727.040 0.000 730.580 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 714.020 0.000 717.560 1.120 ;
  LAYER metal4 ;
  RECT 714.020 0.000 717.560 1.120 ;
  LAYER metal3 ;
  RECT 714.020 0.000 717.560 1.120 ;
  LAYER metal2 ;
  RECT 714.020 0.000 717.560 1.120 ;
  LAYER metal1 ;
  RECT 714.020 0.000 717.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 700.380 0.000 703.920 1.120 ;
  LAYER metal4 ;
  RECT 700.380 0.000 703.920 1.120 ;
  LAYER metal3 ;
  RECT 700.380 0.000 703.920 1.120 ;
  LAYER metal2 ;
  RECT 700.380 0.000 703.920 1.120 ;
  LAYER metal1 ;
  RECT 700.380 0.000 703.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 686.740 0.000 690.280 1.120 ;
  LAYER metal4 ;
  RECT 686.740 0.000 690.280 1.120 ;
  LAYER metal3 ;
  RECT 686.740 0.000 690.280 1.120 ;
  LAYER metal2 ;
  RECT 686.740 0.000 690.280 1.120 ;
  LAYER metal1 ;
  RECT 686.740 0.000 690.280 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 619.780 0.000 623.320 1.120 ;
  LAYER metal4 ;
  RECT 619.780 0.000 623.320 1.120 ;
  LAYER metal3 ;
  RECT 619.780 0.000 623.320 1.120 ;
  LAYER metal2 ;
  RECT 619.780 0.000 623.320 1.120 ;
  LAYER metal1 ;
  RECT 619.780 0.000 623.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 606.140 0.000 609.680 1.120 ;
  LAYER metal4 ;
  RECT 606.140 0.000 609.680 1.120 ;
  LAYER metal3 ;
  RECT 606.140 0.000 609.680 1.120 ;
  LAYER metal2 ;
  RECT 606.140 0.000 609.680 1.120 ;
  LAYER metal1 ;
  RECT 606.140 0.000 609.680 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 593.120 0.000 596.660 1.120 ;
  LAYER metal4 ;
  RECT 593.120 0.000 596.660 1.120 ;
  LAYER metal3 ;
  RECT 593.120 0.000 596.660 1.120 ;
  LAYER metal2 ;
  RECT 593.120 0.000 596.660 1.120 ;
  LAYER metal1 ;
  RECT 593.120 0.000 596.660 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 579.480 0.000 583.020 1.120 ;
  LAYER metal4 ;
  RECT 579.480 0.000 583.020 1.120 ;
  LAYER metal3 ;
  RECT 579.480 0.000 583.020 1.120 ;
  LAYER metal2 ;
  RECT 579.480 0.000 583.020 1.120 ;
  LAYER metal1 ;
  RECT 579.480 0.000 583.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 565.840 0.000 569.380 1.120 ;
  LAYER metal4 ;
  RECT 565.840 0.000 569.380 1.120 ;
  LAYER metal3 ;
  RECT 565.840 0.000 569.380 1.120 ;
  LAYER metal2 ;
  RECT 565.840 0.000 569.380 1.120 ;
  LAYER metal1 ;
  RECT 565.840 0.000 569.380 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 552.820 0.000 556.360 1.120 ;
  LAYER metal4 ;
  RECT 552.820 0.000 556.360 1.120 ;
  LAYER metal3 ;
  RECT 552.820 0.000 556.360 1.120 ;
  LAYER metal2 ;
  RECT 552.820 0.000 556.360 1.120 ;
  LAYER metal1 ;
  RECT 552.820 0.000 556.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 485.240 0.000 488.780 1.120 ;
  LAYER metal4 ;
  RECT 485.240 0.000 488.780 1.120 ;
  LAYER metal3 ;
  RECT 485.240 0.000 488.780 1.120 ;
  LAYER metal2 ;
  RECT 485.240 0.000 488.780 1.120 ;
  LAYER metal1 ;
  RECT 485.240 0.000 488.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 471.600 0.000 475.140 1.120 ;
  LAYER metal4 ;
  RECT 471.600 0.000 475.140 1.120 ;
  LAYER metal3 ;
  RECT 471.600 0.000 475.140 1.120 ;
  LAYER metal2 ;
  RECT 471.600 0.000 475.140 1.120 ;
  LAYER metal1 ;
  RECT 471.600 0.000 475.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 458.580 0.000 462.120 1.120 ;
  LAYER metal4 ;
  RECT 458.580 0.000 462.120 1.120 ;
  LAYER metal3 ;
  RECT 458.580 0.000 462.120 1.120 ;
  LAYER metal2 ;
  RECT 458.580 0.000 462.120 1.120 ;
  LAYER metal1 ;
  RECT 458.580 0.000 462.120 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 444.940 0.000 448.480 1.120 ;
  LAYER metal4 ;
  RECT 444.940 0.000 448.480 1.120 ;
  LAYER metal3 ;
  RECT 444.940 0.000 448.480 1.120 ;
  LAYER metal2 ;
  RECT 444.940 0.000 448.480 1.120 ;
  LAYER metal1 ;
  RECT 444.940 0.000 448.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 431.300 0.000 434.840 1.120 ;
  LAYER metal4 ;
  RECT 431.300 0.000 434.840 1.120 ;
  LAYER metal3 ;
  RECT 431.300 0.000 434.840 1.120 ;
  LAYER metal2 ;
  RECT 431.300 0.000 434.840 1.120 ;
  LAYER metal1 ;
  RECT 431.300 0.000 434.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 418.280 0.000 421.820 1.120 ;
  LAYER metal4 ;
  RECT 418.280 0.000 421.820 1.120 ;
  LAYER metal3 ;
  RECT 418.280 0.000 421.820 1.120 ;
  LAYER metal2 ;
  RECT 418.280 0.000 421.820 1.120 ;
  LAYER metal1 ;
  RECT 418.280 0.000 421.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 350.700 0.000 354.240 1.120 ;
  LAYER metal4 ;
  RECT 350.700 0.000 354.240 1.120 ;
  LAYER metal3 ;
  RECT 350.700 0.000 354.240 1.120 ;
  LAYER metal2 ;
  RECT 350.700 0.000 354.240 1.120 ;
  LAYER metal1 ;
  RECT 350.700 0.000 354.240 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 337.680 0.000 341.220 1.120 ;
  LAYER metal4 ;
  RECT 337.680 0.000 341.220 1.120 ;
  LAYER metal3 ;
  RECT 337.680 0.000 341.220 1.120 ;
  LAYER metal2 ;
  RECT 337.680 0.000 341.220 1.120 ;
  LAYER metal1 ;
  RECT 337.680 0.000 341.220 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 324.040 0.000 327.580 1.120 ;
  LAYER metal4 ;
  RECT 324.040 0.000 327.580 1.120 ;
  LAYER metal3 ;
  RECT 324.040 0.000 327.580 1.120 ;
  LAYER metal2 ;
  RECT 324.040 0.000 327.580 1.120 ;
  LAYER metal1 ;
  RECT 324.040 0.000 327.580 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 310.400 0.000 313.940 1.120 ;
  LAYER metal4 ;
  RECT 310.400 0.000 313.940 1.120 ;
  LAYER metal3 ;
  RECT 310.400 0.000 313.940 1.120 ;
  LAYER metal2 ;
  RECT 310.400 0.000 313.940 1.120 ;
  LAYER metal1 ;
  RECT 310.400 0.000 313.940 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 297.380 0.000 300.920 1.120 ;
  LAYER metal4 ;
  RECT 297.380 0.000 300.920 1.120 ;
  LAYER metal3 ;
  RECT 297.380 0.000 300.920 1.120 ;
  LAYER metal2 ;
  RECT 297.380 0.000 300.920 1.120 ;
  LAYER metal1 ;
  RECT 297.380 0.000 300.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 283.740 0.000 287.280 1.120 ;
  LAYER metal4 ;
  RECT 283.740 0.000 287.280 1.120 ;
  LAYER metal3 ;
  RECT 283.740 0.000 287.280 1.120 ;
  LAYER metal2 ;
  RECT 283.740 0.000 287.280 1.120 ;
  LAYER metal1 ;
  RECT 283.740 0.000 287.280 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 216.780 0.000 220.320 1.120 ;
  LAYER metal4 ;
  RECT 216.780 0.000 220.320 1.120 ;
  LAYER metal3 ;
  RECT 216.780 0.000 220.320 1.120 ;
  LAYER metal2 ;
  RECT 216.780 0.000 220.320 1.120 ;
  LAYER metal1 ;
  RECT 216.780 0.000 220.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 203.140 0.000 206.680 1.120 ;
  LAYER metal4 ;
  RECT 203.140 0.000 206.680 1.120 ;
  LAYER metal3 ;
  RECT 203.140 0.000 206.680 1.120 ;
  LAYER metal2 ;
  RECT 203.140 0.000 206.680 1.120 ;
  LAYER metal1 ;
  RECT 203.140 0.000 206.680 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 189.500 0.000 193.040 1.120 ;
  LAYER metal4 ;
  RECT 189.500 0.000 193.040 1.120 ;
  LAYER metal3 ;
  RECT 189.500 0.000 193.040 1.120 ;
  LAYER metal2 ;
  RECT 189.500 0.000 193.040 1.120 ;
  LAYER metal1 ;
  RECT 189.500 0.000 193.040 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 176.480 0.000 180.020 1.120 ;
  LAYER metal4 ;
  RECT 176.480 0.000 180.020 1.120 ;
  LAYER metal3 ;
  RECT 176.480 0.000 180.020 1.120 ;
  LAYER metal2 ;
  RECT 176.480 0.000 180.020 1.120 ;
  LAYER metal1 ;
  RECT 176.480 0.000 180.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 162.840 0.000 166.380 1.120 ;
  LAYER metal4 ;
  RECT 162.840 0.000 166.380 1.120 ;
  LAYER metal3 ;
  RECT 162.840 0.000 166.380 1.120 ;
  LAYER metal2 ;
  RECT 162.840 0.000 166.380 1.120 ;
  LAYER metal1 ;
  RECT 162.840 0.000 166.380 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 149.200 0.000 152.740 1.120 ;
  LAYER metal4 ;
  RECT 149.200 0.000 152.740 1.120 ;
  LAYER metal3 ;
  RECT 149.200 0.000 152.740 1.120 ;
  LAYER metal2 ;
  RECT 149.200 0.000 152.740 1.120 ;
  LAYER metal1 ;
  RECT 149.200 0.000 152.740 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 82.240 0.000 85.780 1.120 ;
  LAYER metal4 ;
  RECT 82.240 0.000 85.780 1.120 ;
  LAYER metal3 ;
  RECT 82.240 0.000 85.780 1.120 ;
  LAYER metal2 ;
  RECT 82.240 0.000 85.780 1.120 ;
  LAYER metal1 ;
  RECT 82.240 0.000 85.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 68.600 0.000 72.140 1.120 ;
  LAYER metal4 ;
  RECT 68.600 0.000 72.140 1.120 ;
  LAYER metal3 ;
  RECT 68.600 0.000 72.140 1.120 ;
  LAYER metal2 ;
  RECT 68.600 0.000 72.140 1.120 ;
  LAYER metal1 ;
  RECT 68.600 0.000 72.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 54.960 0.000 58.500 1.120 ;
  LAYER metal4 ;
  RECT 54.960 0.000 58.500 1.120 ;
  LAYER metal3 ;
  RECT 54.960 0.000 58.500 1.120 ;
  LAYER metal2 ;
  RECT 54.960 0.000 58.500 1.120 ;
  LAYER metal1 ;
  RECT 54.960 0.000 58.500 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 41.940 0.000 45.480 1.120 ;
  LAYER metal4 ;
  RECT 41.940 0.000 45.480 1.120 ;
  LAYER metal3 ;
  RECT 41.940 0.000 45.480 1.120 ;
  LAYER metal2 ;
  RECT 41.940 0.000 45.480 1.120 ;
  LAYER metal1 ;
  RECT 41.940 0.000 45.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 28.300 0.000 31.840 1.120 ;
  LAYER metal4 ;
  RECT 28.300 0.000 31.840 1.120 ;
  LAYER metal3 ;
  RECT 28.300 0.000 31.840 1.120 ;
  LAYER metal2 ;
  RECT 28.300 0.000 31.840 1.120 ;
  LAYER metal1 ;
  RECT 28.300 0.000 31.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 14.660 0.000 18.200 1.120 ;
  LAYER metal4 ;
  RECT 14.660 0.000 18.200 1.120 ;
  LAYER metal3 ;
  RECT 14.660 0.000 18.200 1.120 ;
  LAYER metal2 ;
  RECT 14.660 0.000 18.200 1.120 ;
  LAYER metal1 ;
  RECT 14.660 0.000 18.200 1.120 ;
 END
END GND
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal5 ;
  RECT 3570.700 195.780 3571.820 199.020 ;
  LAYER metal4 ;
  RECT 3570.700 195.780 3571.820 199.020 ;
  LAYER metal3 ;
  RECT 3570.700 195.780 3571.820 199.020 ;
  LAYER metal2 ;
  RECT 3570.700 195.780 3571.820 199.020 ;
  LAYER metal1 ;
  RECT 3570.700 195.780 3571.820 199.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.700 187.940 3571.820 191.180 ;
  LAYER metal4 ;
  RECT 3570.700 187.940 3571.820 191.180 ;
  LAYER metal3 ;
  RECT 3570.700 187.940 3571.820 191.180 ;
  LAYER metal2 ;
  RECT 3570.700 187.940 3571.820 191.180 ;
  LAYER metal1 ;
  RECT 3570.700 187.940 3571.820 191.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.700 180.100 3571.820 183.340 ;
  LAYER metal4 ;
  RECT 3570.700 180.100 3571.820 183.340 ;
  LAYER metal3 ;
  RECT 3570.700 180.100 3571.820 183.340 ;
  LAYER metal2 ;
  RECT 3570.700 180.100 3571.820 183.340 ;
  LAYER metal1 ;
  RECT 3570.700 180.100 3571.820 183.340 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.700 172.260 3571.820 175.500 ;
  LAYER metal4 ;
  RECT 3570.700 172.260 3571.820 175.500 ;
  LAYER metal3 ;
  RECT 3570.700 172.260 3571.820 175.500 ;
  LAYER metal2 ;
  RECT 3570.700 172.260 3571.820 175.500 ;
  LAYER metal1 ;
  RECT 3570.700 172.260 3571.820 175.500 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.700 164.420 3571.820 167.660 ;
  LAYER metal4 ;
  RECT 3570.700 164.420 3571.820 167.660 ;
  LAYER metal3 ;
  RECT 3570.700 164.420 3571.820 167.660 ;
  LAYER metal2 ;
  RECT 3570.700 164.420 3571.820 167.660 ;
  LAYER metal1 ;
  RECT 3570.700 164.420 3571.820 167.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.700 125.220 3571.820 128.460 ;
  LAYER metal4 ;
  RECT 3570.700 125.220 3571.820 128.460 ;
  LAYER metal3 ;
  RECT 3570.700 125.220 3571.820 128.460 ;
  LAYER metal2 ;
  RECT 3570.700 125.220 3571.820 128.460 ;
  LAYER metal1 ;
  RECT 3570.700 125.220 3571.820 128.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.700 117.380 3571.820 120.620 ;
  LAYER metal4 ;
  RECT 3570.700 117.380 3571.820 120.620 ;
  LAYER metal3 ;
  RECT 3570.700 117.380 3571.820 120.620 ;
  LAYER metal2 ;
  RECT 3570.700 117.380 3571.820 120.620 ;
  LAYER metal1 ;
  RECT 3570.700 117.380 3571.820 120.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.700 109.540 3571.820 112.780 ;
  LAYER metal4 ;
  RECT 3570.700 109.540 3571.820 112.780 ;
  LAYER metal3 ;
  RECT 3570.700 109.540 3571.820 112.780 ;
  LAYER metal2 ;
  RECT 3570.700 109.540 3571.820 112.780 ;
  LAYER metal1 ;
  RECT 3570.700 109.540 3571.820 112.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.700 101.700 3571.820 104.940 ;
  LAYER metal4 ;
  RECT 3570.700 101.700 3571.820 104.940 ;
  LAYER metal3 ;
  RECT 3570.700 101.700 3571.820 104.940 ;
  LAYER metal2 ;
  RECT 3570.700 101.700 3571.820 104.940 ;
  LAYER metal1 ;
  RECT 3570.700 101.700 3571.820 104.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.700 93.860 3571.820 97.100 ;
  LAYER metal4 ;
  RECT 3570.700 93.860 3571.820 97.100 ;
  LAYER metal3 ;
  RECT 3570.700 93.860 3571.820 97.100 ;
  LAYER metal2 ;
  RECT 3570.700 93.860 3571.820 97.100 ;
  LAYER metal1 ;
  RECT 3570.700 93.860 3571.820 97.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.700 86.020 3571.820 89.260 ;
  LAYER metal4 ;
  RECT 3570.700 86.020 3571.820 89.260 ;
  LAYER metal3 ;
  RECT 3570.700 86.020 3571.820 89.260 ;
  LAYER metal2 ;
  RECT 3570.700 86.020 3571.820 89.260 ;
  LAYER metal1 ;
  RECT 3570.700 86.020 3571.820 89.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.700 46.820 3571.820 50.060 ;
  LAYER metal4 ;
  RECT 3570.700 46.820 3571.820 50.060 ;
  LAYER metal3 ;
  RECT 3570.700 46.820 3571.820 50.060 ;
  LAYER metal2 ;
  RECT 3570.700 46.820 3571.820 50.060 ;
  LAYER metal1 ;
  RECT 3570.700 46.820 3571.820 50.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.700 38.980 3571.820 42.220 ;
  LAYER metal4 ;
  RECT 3570.700 38.980 3571.820 42.220 ;
  LAYER metal3 ;
  RECT 3570.700 38.980 3571.820 42.220 ;
  LAYER metal2 ;
  RECT 3570.700 38.980 3571.820 42.220 ;
  LAYER metal1 ;
  RECT 3570.700 38.980 3571.820 42.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.700 31.140 3571.820 34.380 ;
  LAYER metal4 ;
  RECT 3570.700 31.140 3571.820 34.380 ;
  LAYER metal3 ;
  RECT 3570.700 31.140 3571.820 34.380 ;
  LAYER metal2 ;
  RECT 3570.700 31.140 3571.820 34.380 ;
  LAYER metal1 ;
  RECT 3570.700 31.140 3571.820 34.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.700 23.300 3571.820 26.540 ;
  LAYER metal4 ;
  RECT 3570.700 23.300 3571.820 26.540 ;
  LAYER metal3 ;
  RECT 3570.700 23.300 3571.820 26.540 ;
  LAYER metal2 ;
  RECT 3570.700 23.300 3571.820 26.540 ;
  LAYER metal1 ;
  RECT 3570.700 23.300 3571.820 26.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.700 15.460 3571.820 18.700 ;
  LAYER metal4 ;
  RECT 3570.700 15.460 3571.820 18.700 ;
  LAYER metal3 ;
  RECT 3570.700 15.460 3571.820 18.700 ;
  LAYER metal2 ;
  RECT 3570.700 15.460 3571.820 18.700 ;
  LAYER metal1 ;
  RECT 3570.700 15.460 3571.820 18.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3570.700 7.620 3571.820 10.860 ;
  LAYER metal4 ;
  RECT 3570.700 7.620 3571.820 10.860 ;
  LAYER metal3 ;
  RECT 3570.700 7.620 3571.820 10.860 ;
  LAYER metal2 ;
  RECT 3570.700 7.620 3571.820 10.860 ;
  LAYER metal1 ;
  RECT 3570.700 7.620 3571.820 10.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 195.780 1.120 199.020 ;
  LAYER metal4 ;
  RECT 0.000 195.780 1.120 199.020 ;
  LAYER metal3 ;
  RECT 0.000 195.780 1.120 199.020 ;
  LAYER metal2 ;
  RECT 0.000 195.780 1.120 199.020 ;
  LAYER metal1 ;
  RECT 0.000 195.780 1.120 199.020 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 187.940 1.120 191.180 ;
  LAYER metal4 ;
  RECT 0.000 187.940 1.120 191.180 ;
  LAYER metal3 ;
  RECT 0.000 187.940 1.120 191.180 ;
  LAYER metal2 ;
  RECT 0.000 187.940 1.120 191.180 ;
  LAYER metal1 ;
  RECT 0.000 187.940 1.120 191.180 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 180.100 1.120 183.340 ;
  LAYER metal4 ;
  RECT 0.000 180.100 1.120 183.340 ;
  LAYER metal3 ;
  RECT 0.000 180.100 1.120 183.340 ;
  LAYER metal2 ;
  RECT 0.000 180.100 1.120 183.340 ;
  LAYER metal1 ;
  RECT 0.000 180.100 1.120 183.340 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 172.260 1.120 175.500 ;
  LAYER metal4 ;
  RECT 0.000 172.260 1.120 175.500 ;
  LAYER metal3 ;
  RECT 0.000 172.260 1.120 175.500 ;
  LAYER metal2 ;
  RECT 0.000 172.260 1.120 175.500 ;
  LAYER metal1 ;
  RECT 0.000 172.260 1.120 175.500 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 164.420 1.120 167.660 ;
  LAYER metal4 ;
  RECT 0.000 164.420 1.120 167.660 ;
  LAYER metal3 ;
  RECT 0.000 164.420 1.120 167.660 ;
  LAYER metal2 ;
  RECT 0.000 164.420 1.120 167.660 ;
  LAYER metal1 ;
  RECT 0.000 164.420 1.120 167.660 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 125.220 1.120 128.460 ;
  LAYER metal4 ;
  RECT 0.000 125.220 1.120 128.460 ;
  LAYER metal3 ;
  RECT 0.000 125.220 1.120 128.460 ;
  LAYER metal2 ;
  RECT 0.000 125.220 1.120 128.460 ;
  LAYER metal1 ;
  RECT 0.000 125.220 1.120 128.460 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 117.380 1.120 120.620 ;
  LAYER metal4 ;
  RECT 0.000 117.380 1.120 120.620 ;
  LAYER metal3 ;
  RECT 0.000 117.380 1.120 120.620 ;
  LAYER metal2 ;
  RECT 0.000 117.380 1.120 120.620 ;
  LAYER metal1 ;
  RECT 0.000 117.380 1.120 120.620 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 109.540 1.120 112.780 ;
  LAYER metal4 ;
  RECT 0.000 109.540 1.120 112.780 ;
  LAYER metal3 ;
  RECT 0.000 109.540 1.120 112.780 ;
  LAYER metal2 ;
  RECT 0.000 109.540 1.120 112.780 ;
  LAYER metal1 ;
  RECT 0.000 109.540 1.120 112.780 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 101.700 1.120 104.940 ;
  LAYER metal4 ;
  RECT 0.000 101.700 1.120 104.940 ;
  LAYER metal3 ;
  RECT 0.000 101.700 1.120 104.940 ;
  LAYER metal2 ;
  RECT 0.000 101.700 1.120 104.940 ;
  LAYER metal1 ;
  RECT 0.000 101.700 1.120 104.940 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 93.860 1.120 97.100 ;
  LAYER metal4 ;
  RECT 0.000 93.860 1.120 97.100 ;
  LAYER metal3 ;
  RECT 0.000 93.860 1.120 97.100 ;
  LAYER metal2 ;
  RECT 0.000 93.860 1.120 97.100 ;
  LAYER metal1 ;
  RECT 0.000 93.860 1.120 97.100 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 86.020 1.120 89.260 ;
  LAYER metal4 ;
  RECT 0.000 86.020 1.120 89.260 ;
  LAYER metal3 ;
  RECT 0.000 86.020 1.120 89.260 ;
  LAYER metal2 ;
  RECT 0.000 86.020 1.120 89.260 ;
  LAYER metal1 ;
  RECT 0.000 86.020 1.120 89.260 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 46.820 1.120 50.060 ;
  LAYER metal4 ;
  RECT 0.000 46.820 1.120 50.060 ;
  LAYER metal3 ;
  RECT 0.000 46.820 1.120 50.060 ;
  LAYER metal2 ;
  RECT 0.000 46.820 1.120 50.060 ;
  LAYER metal1 ;
  RECT 0.000 46.820 1.120 50.060 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 38.980 1.120 42.220 ;
  LAYER metal4 ;
  RECT 0.000 38.980 1.120 42.220 ;
  LAYER metal3 ;
  RECT 0.000 38.980 1.120 42.220 ;
  LAYER metal2 ;
  RECT 0.000 38.980 1.120 42.220 ;
  LAYER metal1 ;
  RECT 0.000 38.980 1.120 42.220 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 31.140 1.120 34.380 ;
  LAYER metal4 ;
  RECT 0.000 31.140 1.120 34.380 ;
  LAYER metal3 ;
  RECT 0.000 31.140 1.120 34.380 ;
  LAYER metal2 ;
  RECT 0.000 31.140 1.120 34.380 ;
  LAYER metal1 ;
  RECT 0.000 31.140 1.120 34.380 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 23.300 1.120 26.540 ;
  LAYER metal4 ;
  RECT 0.000 23.300 1.120 26.540 ;
  LAYER metal3 ;
  RECT 0.000 23.300 1.120 26.540 ;
  LAYER metal2 ;
  RECT 0.000 23.300 1.120 26.540 ;
  LAYER metal1 ;
  RECT 0.000 23.300 1.120 26.540 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 15.460 1.120 18.700 ;
  LAYER metal4 ;
  RECT 0.000 15.460 1.120 18.700 ;
  LAYER metal3 ;
  RECT 0.000 15.460 1.120 18.700 ;
  LAYER metal2 ;
  RECT 0.000 15.460 1.120 18.700 ;
  LAYER metal1 ;
  RECT 0.000 15.460 1.120 18.700 ;
 END
 PORT
  LAYER metal5 ;
  RECT 0.000 7.620 1.120 10.860 ;
  LAYER metal4 ;
  RECT 0.000 7.620 1.120 10.860 ;
  LAYER metal3 ;
  RECT 0.000 7.620 1.120 10.860 ;
  LAYER metal2 ;
  RECT 0.000 7.620 1.120 10.860 ;
  LAYER metal1 ;
  RECT 0.000 7.620 1.120 10.860 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3559.820 208.880 3563.360 210.000 ;
  LAYER metal4 ;
  RECT 3559.820 208.880 3563.360 210.000 ;
  LAYER metal3 ;
  RECT 3559.820 208.880 3563.360 210.000 ;
  LAYER metal2 ;
  RECT 3559.820 208.880 3563.360 210.000 ;
  LAYER metal1 ;
  RECT 3559.820 208.880 3563.360 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3551.140 208.880 3554.680 210.000 ;
  LAYER metal4 ;
  RECT 3551.140 208.880 3554.680 210.000 ;
  LAYER metal3 ;
  RECT 3551.140 208.880 3554.680 210.000 ;
  LAYER metal2 ;
  RECT 3551.140 208.880 3554.680 210.000 ;
  LAYER metal1 ;
  RECT 3551.140 208.880 3554.680 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3537.500 208.880 3541.040 210.000 ;
  LAYER metal4 ;
  RECT 3537.500 208.880 3541.040 210.000 ;
  LAYER metal3 ;
  RECT 3537.500 208.880 3541.040 210.000 ;
  LAYER metal2 ;
  RECT 3537.500 208.880 3541.040 210.000 ;
  LAYER metal1 ;
  RECT 3537.500 208.880 3541.040 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3524.480 208.880 3528.020 210.000 ;
  LAYER metal4 ;
  RECT 3524.480 208.880 3528.020 210.000 ;
  LAYER metal3 ;
  RECT 3524.480 208.880 3528.020 210.000 ;
  LAYER metal2 ;
  RECT 3524.480 208.880 3528.020 210.000 ;
  LAYER metal1 ;
  RECT 3524.480 208.880 3528.020 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3456.900 208.880 3460.440 210.000 ;
  LAYER metal4 ;
  RECT 3456.900 208.880 3460.440 210.000 ;
  LAYER metal3 ;
  RECT 3456.900 208.880 3460.440 210.000 ;
  LAYER metal2 ;
  RECT 3456.900 208.880 3460.440 210.000 ;
  LAYER metal1 ;
  RECT 3456.900 208.880 3460.440 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3443.260 208.880 3446.800 210.000 ;
  LAYER metal4 ;
  RECT 3443.260 208.880 3446.800 210.000 ;
  LAYER metal3 ;
  RECT 3443.260 208.880 3446.800 210.000 ;
  LAYER metal2 ;
  RECT 3443.260 208.880 3446.800 210.000 ;
  LAYER metal1 ;
  RECT 3443.260 208.880 3446.800 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3430.240 208.880 3433.780 210.000 ;
  LAYER metal4 ;
  RECT 3430.240 208.880 3433.780 210.000 ;
  LAYER metal3 ;
  RECT 3430.240 208.880 3433.780 210.000 ;
  LAYER metal2 ;
  RECT 3430.240 208.880 3433.780 210.000 ;
  LAYER metal1 ;
  RECT 3430.240 208.880 3433.780 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3416.600 208.880 3420.140 210.000 ;
  LAYER metal4 ;
  RECT 3416.600 208.880 3420.140 210.000 ;
  LAYER metal3 ;
  RECT 3416.600 208.880 3420.140 210.000 ;
  LAYER metal2 ;
  RECT 3416.600 208.880 3420.140 210.000 ;
  LAYER metal1 ;
  RECT 3416.600 208.880 3420.140 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3402.960 208.880 3406.500 210.000 ;
  LAYER metal4 ;
  RECT 3402.960 208.880 3406.500 210.000 ;
  LAYER metal3 ;
  RECT 3402.960 208.880 3406.500 210.000 ;
  LAYER metal2 ;
  RECT 3402.960 208.880 3406.500 210.000 ;
  LAYER metal1 ;
  RECT 3402.960 208.880 3406.500 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3389.940 208.880 3393.480 210.000 ;
  LAYER metal4 ;
  RECT 3389.940 208.880 3393.480 210.000 ;
  LAYER metal3 ;
  RECT 3389.940 208.880 3393.480 210.000 ;
  LAYER metal2 ;
  RECT 3389.940 208.880 3393.480 210.000 ;
  LAYER metal1 ;
  RECT 3389.940 208.880 3393.480 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3322.360 208.880 3325.900 210.000 ;
  LAYER metal4 ;
  RECT 3322.360 208.880 3325.900 210.000 ;
  LAYER metal3 ;
  RECT 3322.360 208.880 3325.900 210.000 ;
  LAYER metal2 ;
  RECT 3322.360 208.880 3325.900 210.000 ;
  LAYER metal1 ;
  RECT 3322.360 208.880 3325.900 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3309.340 208.880 3312.880 210.000 ;
  LAYER metal4 ;
  RECT 3309.340 208.880 3312.880 210.000 ;
  LAYER metal3 ;
  RECT 3309.340 208.880 3312.880 210.000 ;
  LAYER metal2 ;
  RECT 3309.340 208.880 3312.880 210.000 ;
  LAYER metal1 ;
  RECT 3309.340 208.880 3312.880 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3295.700 208.880 3299.240 210.000 ;
  LAYER metal4 ;
  RECT 3295.700 208.880 3299.240 210.000 ;
  LAYER metal3 ;
  RECT 3295.700 208.880 3299.240 210.000 ;
  LAYER metal2 ;
  RECT 3295.700 208.880 3299.240 210.000 ;
  LAYER metal1 ;
  RECT 3295.700 208.880 3299.240 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3282.060 208.880 3285.600 210.000 ;
  LAYER metal4 ;
  RECT 3282.060 208.880 3285.600 210.000 ;
  LAYER metal3 ;
  RECT 3282.060 208.880 3285.600 210.000 ;
  LAYER metal2 ;
  RECT 3282.060 208.880 3285.600 210.000 ;
  LAYER metal1 ;
  RECT 3282.060 208.880 3285.600 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3269.040 208.880 3272.580 210.000 ;
  LAYER metal4 ;
  RECT 3269.040 208.880 3272.580 210.000 ;
  LAYER metal3 ;
  RECT 3269.040 208.880 3272.580 210.000 ;
  LAYER metal2 ;
  RECT 3269.040 208.880 3272.580 210.000 ;
  LAYER metal1 ;
  RECT 3269.040 208.880 3272.580 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3255.400 208.880 3258.940 210.000 ;
  LAYER metal4 ;
  RECT 3255.400 208.880 3258.940 210.000 ;
  LAYER metal3 ;
  RECT 3255.400 208.880 3258.940 210.000 ;
  LAYER metal2 ;
  RECT 3255.400 208.880 3258.940 210.000 ;
  LAYER metal1 ;
  RECT 3255.400 208.880 3258.940 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3188.440 208.880 3191.980 210.000 ;
  LAYER metal4 ;
  RECT 3188.440 208.880 3191.980 210.000 ;
  LAYER metal3 ;
  RECT 3188.440 208.880 3191.980 210.000 ;
  LAYER metal2 ;
  RECT 3188.440 208.880 3191.980 210.000 ;
  LAYER metal1 ;
  RECT 3188.440 208.880 3191.980 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3174.800 208.880 3178.340 210.000 ;
  LAYER metal4 ;
  RECT 3174.800 208.880 3178.340 210.000 ;
  LAYER metal3 ;
  RECT 3174.800 208.880 3178.340 210.000 ;
  LAYER metal2 ;
  RECT 3174.800 208.880 3178.340 210.000 ;
  LAYER metal1 ;
  RECT 3174.800 208.880 3178.340 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3161.160 208.880 3164.700 210.000 ;
  LAYER metal4 ;
  RECT 3161.160 208.880 3164.700 210.000 ;
  LAYER metal3 ;
  RECT 3161.160 208.880 3164.700 210.000 ;
  LAYER metal2 ;
  RECT 3161.160 208.880 3164.700 210.000 ;
  LAYER metal1 ;
  RECT 3161.160 208.880 3164.700 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3148.140 208.880 3151.680 210.000 ;
  LAYER metal4 ;
  RECT 3148.140 208.880 3151.680 210.000 ;
  LAYER metal3 ;
  RECT 3148.140 208.880 3151.680 210.000 ;
  LAYER metal2 ;
  RECT 3148.140 208.880 3151.680 210.000 ;
  LAYER metal1 ;
  RECT 3148.140 208.880 3151.680 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3134.500 208.880 3138.040 210.000 ;
  LAYER metal4 ;
  RECT 3134.500 208.880 3138.040 210.000 ;
  LAYER metal3 ;
  RECT 3134.500 208.880 3138.040 210.000 ;
  LAYER metal2 ;
  RECT 3134.500 208.880 3138.040 210.000 ;
  LAYER metal1 ;
  RECT 3134.500 208.880 3138.040 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3120.860 208.880 3124.400 210.000 ;
  LAYER metal4 ;
  RECT 3120.860 208.880 3124.400 210.000 ;
  LAYER metal3 ;
  RECT 3120.860 208.880 3124.400 210.000 ;
  LAYER metal2 ;
  RECT 3120.860 208.880 3124.400 210.000 ;
  LAYER metal1 ;
  RECT 3120.860 208.880 3124.400 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3053.900 208.880 3057.440 210.000 ;
  LAYER metal4 ;
  RECT 3053.900 208.880 3057.440 210.000 ;
  LAYER metal3 ;
  RECT 3053.900 208.880 3057.440 210.000 ;
  LAYER metal2 ;
  RECT 3053.900 208.880 3057.440 210.000 ;
  LAYER metal1 ;
  RECT 3053.900 208.880 3057.440 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3040.260 208.880 3043.800 210.000 ;
  LAYER metal4 ;
  RECT 3040.260 208.880 3043.800 210.000 ;
  LAYER metal3 ;
  RECT 3040.260 208.880 3043.800 210.000 ;
  LAYER metal2 ;
  RECT 3040.260 208.880 3043.800 210.000 ;
  LAYER metal1 ;
  RECT 3040.260 208.880 3043.800 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3026.620 208.880 3030.160 210.000 ;
  LAYER metal4 ;
  RECT 3026.620 208.880 3030.160 210.000 ;
  LAYER metal3 ;
  RECT 3026.620 208.880 3030.160 210.000 ;
  LAYER metal2 ;
  RECT 3026.620 208.880 3030.160 210.000 ;
  LAYER metal1 ;
  RECT 3026.620 208.880 3030.160 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3013.600 208.880 3017.140 210.000 ;
  LAYER metal4 ;
  RECT 3013.600 208.880 3017.140 210.000 ;
  LAYER metal3 ;
  RECT 3013.600 208.880 3017.140 210.000 ;
  LAYER metal2 ;
  RECT 3013.600 208.880 3017.140 210.000 ;
  LAYER metal1 ;
  RECT 3013.600 208.880 3017.140 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2999.960 208.880 3003.500 210.000 ;
  LAYER metal4 ;
  RECT 2999.960 208.880 3003.500 210.000 ;
  LAYER metal3 ;
  RECT 2999.960 208.880 3003.500 210.000 ;
  LAYER metal2 ;
  RECT 2999.960 208.880 3003.500 210.000 ;
  LAYER metal1 ;
  RECT 2999.960 208.880 3003.500 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2986.320 208.880 2989.860 210.000 ;
  LAYER metal4 ;
  RECT 2986.320 208.880 2989.860 210.000 ;
  LAYER metal3 ;
  RECT 2986.320 208.880 2989.860 210.000 ;
  LAYER metal2 ;
  RECT 2986.320 208.880 2989.860 210.000 ;
  LAYER metal1 ;
  RECT 2986.320 208.880 2989.860 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2919.360 208.880 2922.900 210.000 ;
  LAYER metal4 ;
  RECT 2919.360 208.880 2922.900 210.000 ;
  LAYER metal3 ;
  RECT 2919.360 208.880 2922.900 210.000 ;
  LAYER metal2 ;
  RECT 2919.360 208.880 2922.900 210.000 ;
  LAYER metal1 ;
  RECT 2919.360 208.880 2922.900 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2905.720 208.880 2909.260 210.000 ;
  LAYER metal4 ;
  RECT 2905.720 208.880 2909.260 210.000 ;
  LAYER metal3 ;
  RECT 2905.720 208.880 2909.260 210.000 ;
  LAYER metal2 ;
  RECT 2905.720 208.880 2909.260 210.000 ;
  LAYER metal1 ;
  RECT 2905.720 208.880 2909.260 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2892.700 208.880 2896.240 210.000 ;
  LAYER metal4 ;
  RECT 2892.700 208.880 2896.240 210.000 ;
  LAYER metal3 ;
  RECT 2892.700 208.880 2896.240 210.000 ;
  LAYER metal2 ;
  RECT 2892.700 208.880 2896.240 210.000 ;
  LAYER metal1 ;
  RECT 2892.700 208.880 2896.240 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2879.060 208.880 2882.600 210.000 ;
  LAYER metal4 ;
  RECT 2879.060 208.880 2882.600 210.000 ;
  LAYER metal3 ;
  RECT 2879.060 208.880 2882.600 210.000 ;
  LAYER metal2 ;
  RECT 2879.060 208.880 2882.600 210.000 ;
  LAYER metal1 ;
  RECT 2879.060 208.880 2882.600 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2865.420 208.880 2868.960 210.000 ;
  LAYER metal4 ;
  RECT 2865.420 208.880 2868.960 210.000 ;
  LAYER metal3 ;
  RECT 2865.420 208.880 2868.960 210.000 ;
  LAYER metal2 ;
  RECT 2865.420 208.880 2868.960 210.000 ;
  LAYER metal1 ;
  RECT 2865.420 208.880 2868.960 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2852.400 208.880 2855.940 210.000 ;
  LAYER metal4 ;
  RECT 2852.400 208.880 2855.940 210.000 ;
  LAYER metal3 ;
  RECT 2852.400 208.880 2855.940 210.000 ;
  LAYER metal2 ;
  RECT 2852.400 208.880 2855.940 210.000 ;
  LAYER metal1 ;
  RECT 2852.400 208.880 2855.940 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2784.820 208.880 2788.360 210.000 ;
  LAYER metal4 ;
  RECT 2784.820 208.880 2788.360 210.000 ;
  LAYER metal3 ;
  RECT 2784.820 208.880 2788.360 210.000 ;
  LAYER metal2 ;
  RECT 2784.820 208.880 2788.360 210.000 ;
  LAYER metal1 ;
  RECT 2784.820 208.880 2788.360 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2771.800 208.880 2775.340 210.000 ;
  LAYER metal4 ;
  RECT 2771.800 208.880 2775.340 210.000 ;
  LAYER metal3 ;
  RECT 2771.800 208.880 2775.340 210.000 ;
  LAYER metal2 ;
  RECT 2771.800 208.880 2775.340 210.000 ;
  LAYER metal1 ;
  RECT 2771.800 208.880 2775.340 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2758.160 208.880 2761.700 210.000 ;
  LAYER metal4 ;
  RECT 2758.160 208.880 2761.700 210.000 ;
  LAYER metal3 ;
  RECT 2758.160 208.880 2761.700 210.000 ;
  LAYER metal2 ;
  RECT 2758.160 208.880 2761.700 210.000 ;
  LAYER metal1 ;
  RECT 2758.160 208.880 2761.700 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2744.520 208.880 2748.060 210.000 ;
  LAYER metal4 ;
  RECT 2744.520 208.880 2748.060 210.000 ;
  LAYER metal3 ;
  RECT 2744.520 208.880 2748.060 210.000 ;
  LAYER metal2 ;
  RECT 2744.520 208.880 2748.060 210.000 ;
  LAYER metal1 ;
  RECT 2744.520 208.880 2748.060 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2731.500 208.880 2735.040 210.000 ;
  LAYER metal4 ;
  RECT 2731.500 208.880 2735.040 210.000 ;
  LAYER metal3 ;
  RECT 2731.500 208.880 2735.040 210.000 ;
  LAYER metal2 ;
  RECT 2731.500 208.880 2735.040 210.000 ;
  LAYER metal1 ;
  RECT 2731.500 208.880 2735.040 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2717.860 208.880 2721.400 210.000 ;
  LAYER metal4 ;
  RECT 2717.860 208.880 2721.400 210.000 ;
  LAYER metal3 ;
  RECT 2717.860 208.880 2721.400 210.000 ;
  LAYER metal2 ;
  RECT 2717.860 208.880 2721.400 210.000 ;
  LAYER metal1 ;
  RECT 2717.860 208.880 2721.400 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2650.900 208.880 2654.440 210.000 ;
  LAYER metal4 ;
  RECT 2650.900 208.880 2654.440 210.000 ;
  LAYER metal3 ;
  RECT 2650.900 208.880 2654.440 210.000 ;
  LAYER metal2 ;
  RECT 2650.900 208.880 2654.440 210.000 ;
  LAYER metal1 ;
  RECT 2650.900 208.880 2654.440 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2637.260 208.880 2640.800 210.000 ;
  LAYER metal4 ;
  RECT 2637.260 208.880 2640.800 210.000 ;
  LAYER metal3 ;
  RECT 2637.260 208.880 2640.800 210.000 ;
  LAYER metal2 ;
  RECT 2637.260 208.880 2640.800 210.000 ;
  LAYER metal1 ;
  RECT 2637.260 208.880 2640.800 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2623.620 208.880 2627.160 210.000 ;
  LAYER metal4 ;
  RECT 2623.620 208.880 2627.160 210.000 ;
  LAYER metal3 ;
  RECT 2623.620 208.880 2627.160 210.000 ;
  LAYER metal2 ;
  RECT 2623.620 208.880 2627.160 210.000 ;
  LAYER metal1 ;
  RECT 2623.620 208.880 2627.160 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2609.980 208.880 2613.520 210.000 ;
  LAYER metal4 ;
  RECT 2609.980 208.880 2613.520 210.000 ;
  LAYER metal3 ;
  RECT 2609.980 208.880 2613.520 210.000 ;
  LAYER metal2 ;
  RECT 2609.980 208.880 2613.520 210.000 ;
  LAYER metal1 ;
  RECT 2609.980 208.880 2613.520 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2596.960 208.880 2600.500 210.000 ;
  LAYER metal4 ;
  RECT 2596.960 208.880 2600.500 210.000 ;
  LAYER metal3 ;
  RECT 2596.960 208.880 2600.500 210.000 ;
  LAYER metal2 ;
  RECT 2596.960 208.880 2600.500 210.000 ;
  LAYER metal1 ;
  RECT 2596.960 208.880 2600.500 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2583.320 208.880 2586.860 210.000 ;
  LAYER metal4 ;
  RECT 2583.320 208.880 2586.860 210.000 ;
  LAYER metal3 ;
  RECT 2583.320 208.880 2586.860 210.000 ;
  LAYER metal2 ;
  RECT 2583.320 208.880 2586.860 210.000 ;
  LAYER metal1 ;
  RECT 2583.320 208.880 2586.860 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2516.360 208.880 2519.900 210.000 ;
  LAYER metal4 ;
  RECT 2516.360 208.880 2519.900 210.000 ;
  LAYER metal3 ;
  RECT 2516.360 208.880 2519.900 210.000 ;
  LAYER metal2 ;
  RECT 2516.360 208.880 2519.900 210.000 ;
  LAYER metal1 ;
  RECT 2516.360 208.880 2519.900 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2502.720 208.880 2506.260 210.000 ;
  LAYER metal4 ;
  RECT 2502.720 208.880 2506.260 210.000 ;
  LAYER metal3 ;
  RECT 2502.720 208.880 2506.260 210.000 ;
  LAYER metal2 ;
  RECT 2502.720 208.880 2506.260 210.000 ;
  LAYER metal1 ;
  RECT 2502.720 208.880 2506.260 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2489.080 208.880 2492.620 210.000 ;
  LAYER metal4 ;
  RECT 2489.080 208.880 2492.620 210.000 ;
  LAYER metal3 ;
  RECT 2489.080 208.880 2492.620 210.000 ;
  LAYER metal2 ;
  RECT 2489.080 208.880 2492.620 210.000 ;
  LAYER metal1 ;
  RECT 2489.080 208.880 2492.620 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2476.060 208.880 2479.600 210.000 ;
  LAYER metal4 ;
  RECT 2476.060 208.880 2479.600 210.000 ;
  LAYER metal3 ;
  RECT 2476.060 208.880 2479.600 210.000 ;
  LAYER metal2 ;
  RECT 2476.060 208.880 2479.600 210.000 ;
  LAYER metal1 ;
  RECT 2476.060 208.880 2479.600 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2462.420 208.880 2465.960 210.000 ;
  LAYER metal4 ;
  RECT 2462.420 208.880 2465.960 210.000 ;
  LAYER metal3 ;
  RECT 2462.420 208.880 2465.960 210.000 ;
  LAYER metal2 ;
  RECT 2462.420 208.880 2465.960 210.000 ;
  LAYER metal1 ;
  RECT 2462.420 208.880 2465.960 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2448.780 208.880 2452.320 210.000 ;
  LAYER metal4 ;
  RECT 2448.780 208.880 2452.320 210.000 ;
  LAYER metal3 ;
  RECT 2448.780 208.880 2452.320 210.000 ;
  LAYER metal2 ;
  RECT 2448.780 208.880 2452.320 210.000 ;
  LAYER metal1 ;
  RECT 2448.780 208.880 2452.320 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2381.820 208.880 2385.360 210.000 ;
  LAYER metal4 ;
  RECT 2381.820 208.880 2385.360 210.000 ;
  LAYER metal3 ;
  RECT 2381.820 208.880 2385.360 210.000 ;
  LAYER metal2 ;
  RECT 2381.820 208.880 2385.360 210.000 ;
  LAYER metal1 ;
  RECT 2381.820 208.880 2385.360 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2368.180 208.880 2371.720 210.000 ;
  LAYER metal4 ;
  RECT 2368.180 208.880 2371.720 210.000 ;
  LAYER metal3 ;
  RECT 2368.180 208.880 2371.720 210.000 ;
  LAYER metal2 ;
  RECT 2368.180 208.880 2371.720 210.000 ;
  LAYER metal1 ;
  RECT 2368.180 208.880 2371.720 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2355.160 208.880 2358.700 210.000 ;
  LAYER metal4 ;
  RECT 2355.160 208.880 2358.700 210.000 ;
  LAYER metal3 ;
  RECT 2355.160 208.880 2358.700 210.000 ;
  LAYER metal2 ;
  RECT 2355.160 208.880 2358.700 210.000 ;
  LAYER metal1 ;
  RECT 2355.160 208.880 2358.700 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2341.520 208.880 2345.060 210.000 ;
  LAYER metal4 ;
  RECT 2341.520 208.880 2345.060 210.000 ;
  LAYER metal3 ;
  RECT 2341.520 208.880 2345.060 210.000 ;
  LAYER metal2 ;
  RECT 2341.520 208.880 2345.060 210.000 ;
  LAYER metal1 ;
  RECT 2341.520 208.880 2345.060 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2327.880 208.880 2331.420 210.000 ;
  LAYER metal4 ;
  RECT 2327.880 208.880 2331.420 210.000 ;
  LAYER metal3 ;
  RECT 2327.880 208.880 2331.420 210.000 ;
  LAYER metal2 ;
  RECT 2327.880 208.880 2331.420 210.000 ;
  LAYER metal1 ;
  RECT 2327.880 208.880 2331.420 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2314.860 208.880 2318.400 210.000 ;
  LAYER metal4 ;
  RECT 2314.860 208.880 2318.400 210.000 ;
  LAYER metal3 ;
  RECT 2314.860 208.880 2318.400 210.000 ;
  LAYER metal2 ;
  RECT 2314.860 208.880 2318.400 210.000 ;
  LAYER metal1 ;
  RECT 2314.860 208.880 2318.400 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2247.280 208.880 2250.820 210.000 ;
  LAYER metal4 ;
  RECT 2247.280 208.880 2250.820 210.000 ;
  LAYER metal3 ;
  RECT 2247.280 208.880 2250.820 210.000 ;
  LAYER metal2 ;
  RECT 2247.280 208.880 2250.820 210.000 ;
  LAYER metal1 ;
  RECT 2247.280 208.880 2250.820 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2234.260 208.880 2237.800 210.000 ;
  LAYER metal4 ;
  RECT 2234.260 208.880 2237.800 210.000 ;
  LAYER metal3 ;
  RECT 2234.260 208.880 2237.800 210.000 ;
  LAYER metal2 ;
  RECT 2234.260 208.880 2237.800 210.000 ;
  LAYER metal1 ;
  RECT 2234.260 208.880 2237.800 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2220.620 208.880 2224.160 210.000 ;
  LAYER metal4 ;
  RECT 2220.620 208.880 2224.160 210.000 ;
  LAYER metal3 ;
  RECT 2220.620 208.880 2224.160 210.000 ;
  LAYER metal2 ;
  RECT 2220.620 208.880 2224.160 210.000 ;
  LAYER metal1 ;
  RECT 2220.620 208.880 2224.160 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2206.980 208.880 2210.520 210.000 ;
  LAYER metal4 ;
  RECT 2206.980 208.880 2210.520 210.000 ;
  LAYER metal3 ;
  RECT 2206.980 208.880 2210.520 210.000 ;
  LAYER metal2 ;
  RECT 2206.980 208.880 2210.520 210.000 ;
  LAYER metal1 ;
  RECT 2206.980 208.880 2210.520 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2193.340 208.880 2196.880 210.000 ;
  LAYER metal4 ;
  RECT 2193.340 208.880 2196.880 210.000 ;
  LAYER metal3 ;
  RECT 2193.340 208.880 2196.880 210.000 ;
  LAYER metal2 ;
  RECT 2193.340 208.880 2196.880 210.000 ;
  LAYER metal1 ;
  RECT 2193.340 208.880 2196.880 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2180.320 208.880 2183.860 210.000 ;
  LAYER metal4 ;
  RECT 2180.320 208.880 2183.860 210.000 ;
  LAYER metal3 ;
  RECT 2180.320 208.880 2183.860 210.000 ;
  LAYER metal2 ;
  RECT 2180.320 208.880 2183.860 210.000 ;
  LAYER metal1 ;
  RECT 2180.320 208.880 2183.860 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2112.740 208.880 2116.280 210.000 ;
  LAYER metal4 ;
  RECT 2112.740 208.880 2116.280 210.000 ;
  LAYER metal3 ;
  RECT 2112.740 208.880 2116.280 210.000 ;
  LAYER metal2 ;
  RECT 2112.740 208.880 2116.280 210.000 ;
  LAYER metal1 ;
  RECT 2112.740 208.880 2116.280 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2099.720 208.880 2103.260 210.000 ;
  LAYER metal4 ;
  RECT 2099.720 208.880 2103.260 210.000 ;
  LAYER metal3 ;
  RECT 2099.720 208.880 2103.260 210.000 ;
  LAYER metal2 ;
  RECT 2099.720 208.880 2103.260 210.000 ;
  LAYER metal1 ;
  RECT 2099.720 208.880 2103.260 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2086.080 208.880 2089.620 210.000 ;
  LAYER metal4 ;
  RECT 2086.080 208.880 2089.620 210.000 ;
  LAYER metal3 ;
  RECT 2086.080 208.880 2089.620 210.000 ;
  LAYER metal2 ;
  RECT 2086.080 208.880 2089.620 210.000 ;
  LAYER metal1 ;
  RECT 2086.080 208.880 2089.620 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2072.440 208.880 2075.980 210.000 ;
  LAYER metal4 ;
  RECT 2072.440 208.880 2075.980 210.000 ;
  LAYER metal3 ;
  RECT 2072.440 208.880 2075.980 210.000 ;
  LAYER metal2 ;
  RECT 2072.440 208.880 2075.980 210.000 ;
  LAYER metal1 ;
  RECT 2072.440 208.880 2075.980 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2059.420 208.880 2062.960 210.000 ;
  LAYER metal4 ;
  RECT 2059.420 208.880 2062.960 210.000 ;
  LAYER metal3 ;
  RECT 2059.420 208.880 2062.960 210.000 ;
  LAYER metal2 ;
  RECT 2059.420 208.880 2062.960 210.000 ;
  LAYER metal1 ;
  RECT 2059.420 208.880 2062.960 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2045.780 208.880 2049.320 210.000 ;
  LAYER metal4 ;
  RECT 2045.780 208.880 2049.320 210.000 ;
  LAYER metal3 ;
  RECT 2045.780 208.880 2049.320 210.000 ;
  LAYER metal2 ;
  RECT 2045.780 208.880 2049.320 210.000 ;
  LAYER metal1 ;
  RECT 2045.780 208.880 2049.320 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1978.820 208.880 1982.360 210.000 ;
  LAYER metal4 ;
  RECT 1978.820 208.880 1982.360 210.000 ;
  LAYER metal3 ;
  RECT 1978.820 208.880 1982.360 210.000 ;
  LAYER metal2 ;
  RECT 1978.820 208.880 1982.360 210.000 ;
  LAYER metal1 ;
  RECT 1978.820 208.880 1982.360 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1965.180 208.880 1968.720 210.000 ;
  LAYER metal4 ;
  RECT 1965.180 208.880 1968.720 210.000 ;
  LAYER metal3 ;
  RECT 1965.180 208.880 1968.720 210.000 ;
  LAYER metal2 ;
  RECT 1965.180 208.880 1968.720 210.000 ;
  LAYER metal1 ;
  RECT 1965.180 208.880 1968.720 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1951.540 208.880 1955.080 210.000 ;
  LAYER metal4 ;
  RECT 1951.540 208.880 1955.080 210.000 ;
  LAYER metal3 ;
  RECT 1951.540 208.880 1955.080 210.000 ;
  LAYER metal2 ;
  RECT 1951.540 208.880 1955.080 210.000 ;
  LAYER metal1 ;
  RECT 1951.540 208.880 1955.080 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1938.520 208.880 1942.060 210.000 ;
  LAYER metal4 ;
  RECT 1938.520 208.880 1942.060 210.000 ;
  LAYER metal3 ;
  RECT 1938.520 208.880 1942.060 210.000 ;
  LAYER metal2 ;
  RECT 1938.520 208.880 1942.060 210.000 ;
  LAYER metal1 ;
  RECT 1938.520 208.880 1942.060 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1924.880 208.880 1928.420 210.000 ;
  LAYER metal4 ;
  RECT 1924.880 208.880 1928.420 210.000 ;
  LAYER metal3 ;
  RECT 1924.880 208.880 1928.420 210.000 ;
  LAYER metal2 ;
  RECT 1924.880 208.880 1928.420 210.000 ;
  LAYER metal1 ;
  RECT 1924.880 208.880 1928.420 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1911.240 208.880 1914.780 210.000 ;
  LAYER metal4 ;
  RECT 1911.240 208.880 1914.780 210.000 ;
  LAYER metal3 ;
  RECT 1911.240 208.880 1914.780 210.000 ;
  LAYER metal2 ;
  RECT 1911.240 208.880 1914.780 210.000 ;
  LAYER metal1 ;
  RECT 1911.240 208.880 1914.780 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1844.280 208.880 1847.820 210.000 ;
  LAYER metal4 ;
  RECT 1844.280 208.880 1847.820 210.000 ;
  LAYER metal3 ;
  RECT 1844.280 208.880 1847.820 210.000 ;
  LAYER metal2 ;
  RECT 1844.280 208.880 1847.820 210.000 ;
  LAYER metal1 ;
  RECT 1844.280 208.880 1847.820 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1830.640 208.880 1834.180 210.000 ;
  LAYER metal4 ;
  RECT 1830.640 208.880 1834.180 210.000 ;
  LAYER metal3 ;
  RECT 1830.640 208.880 1834.180 210.000 ;
  LAYER metal2 ;
  RECT 1830.640 208.880 1834.180 210.000 ;
  LAYER metal1 ;
  RECT 1830.640 208.880 1834.180 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1821.960 208.880 1825.500 210.000 ;
  LAYER metal4 ;
  RECT 1821.960 208.880 1825.500 210.000 ;
  LAYER metal3 ;
  RECT 1821.960 208.880 1825.500 210.000 ;
  LAYER metal2 ;
  RECT 1821.960 208.880 1825.500 210.000 ;
  LAYER metal1 ;
  RECT 1821.960 208.880 1825.500 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1808.320 208.880 1811.860 210.000 ;
  LAYER metal4 ;
  RECT 1808.320 208.880 1811.860 210.000 ;
  LAYER metal3 ;
  RECT 1808.320 208.880 1811.860 210.000 ;
  LAYER metal2 ;
  RECT 1808.320 208.880 1811.860 210.000 ;
  LAYER metal1 ;
  RECT 1808.320 208.880 1811.860 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1779.800 208.880 1783.340 210.000 ;
  LAYER metal4 ;
  RECT 1779.800 208.880 1783.340 210.000 ;
  LAYER metal3 ;
  RECT 1779.800 208.880 1783.340 210.000 ;
  LAYER metal2 ;
  RECT 1779.800 208.880 1783.340 210.000 ;
  LAYER metal1 ;
  RECT 1779.800 208.880 1783.340 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1754.380 208.880 1757.920 210.000 ;
  LAYER metal4 ;
  RECT 1754.380 208.880 1757.920 210.000 ;
  LAYER metal3 ;
  RECT 1754.380 208.880 1757.920 210.000 ;
  LAYER metal2 ;
  RECT 1754.380 208.880 1757.920 210.000 ;
  LAYER metal1 ;
  RECT 1754.380 208.880 1757.920 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1685.560 208.880 1689.100 210.000 ;
  LAYER metal4 ;
  RECT 1685.560 208.880 1689.100 210.000 ;
  LAYER metal3 ;
  RECT 1685.560 208.880 1689.100 210.000 ;
  LAYER metal2 ;
  RECT 1685.560 208.880 1689.100 210.000 ;
  LAYER metal1 ;
  RECT 1685.560 208.880 1689.100 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1672.540 208.880 1676.080 210.000 ;
  LAYER metal4 ;
  RECT 1672.540 208.880 1676.080 210.000 ;
  LAYER metal3 ;
  RECT 1672.540 208.880 1676.080 210.000 ;
  LAYER metal2 ;
  RECT 1672.540 208.880 1676.080 210.000 ;
  LAYER metal1 ;
  RECT 1672.540 208.880 1676.080 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1658.900 208.880 1662.440 210.000 ;
  LAYER metal4 ;
  RECT 1658.900 208.880 1662.440 210.000 ;
  LAYER metal3 ;
  RECT 1658.900 208.880 1662.440 210.000 ;
  LAYER metal2 ;
  RECT 1658.900 208.880 1662.440 210.000 ;
  LAYER metal1 ;
  RECT 1658.900 208.880 1662.440 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1645.260 208.880 1648.800 210.000 ;
  LAYER metal4 ;
  RECT 1645.260 208.880 1648.800 210.000 ;
  LAYER metal3 ;
  RECT 1645.260 208.880 1648.800 210.000 ;
  LAYER metal2 ;
  RECT 1645.260 208.880 1648.800 210.000 ;
  LAYER metal1 ;
  RECT 1645.260 208.880 1648.800 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1632.240 208.880 1635.780 210.000 ;
  LAYER metal4 ;
  RECT 1632.240 208.880 1635.780 210.000 ;
  LAYER metal3 ;
  RECT 1632.240 208.880 1635.780 210.000 ;
  LAYER metal2 ;
  RECT 1632.240 208.880 1635.780 210.000 ;
  LAYER metal1 ;
  RECT 1632.240 208.880 1635.780 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1618.600 208.880 1622.140 210.000 ;
  LAYER metal4 ;
  RECT 1618.600 208.880 1622.140 210.000 ;
  LAYER metal3 ;
  RECT 1618.600 208.880 1622.140 210.000 ;
  LAYER metal2 ;
  RECT 1618.600 208.880 1622.140 210.000 ;
  LAYER metal1 ;
  RECT 1618.600 208.880 1622.140 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1551.640 208.880 1555.180 210.000 ;
  LAYER metal4 ;
  RECT 1551.640 208.880 1555.180 210.000 ;
  LAYER metal3 ;
  RECT 1551.640 208.880 1555.180 210.000 ;
  LAYER metal2 ;
  RECT 1551.640 208.880 1555.180 210.000 ;
  LAYER metal1 ;
  RECT 1551.640 208.880 1555.180 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1538.000 208.880 1541.540 210.000 ;
  LAYER metal4 ;
  RECT 1538.000 208.880 1541.540 210.000 ;
  LAYER metal3 ;
  RECT 1538.000 208.880 1541.540 210.000 ;
  LAYER metal2 ;
  RECT 1538.000 208.880 1541.540 210.000 ;
  LAYER metal1 ;
  RECT 1538.000 208.880 1541.540 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1524.360 208.880 1527.900 210.000 ;
  LAYER metal4 ;
  RECT 1524.360 208.880 1527.900 210.000 ;
  LAYER metal3 ;
  RECT 1524.360 208.880 1527.900 210.000 ;
  LAYER metal2 ;
  RECT 1524.360 208.880 1527.900 210.000 ;
  LAYER metal1 ;
  RECT 1524.360 208.880 1527.900 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1511.340 208.880 1514.880 210.000 ;
  LAYER metal4 ;
  RECT 1511.340 208.880 1514.880 210.000 ;
  LAYER metal3 ;
  RECT 1511.340 208.880 1514.880 210.000 ;
  LAYER metal2 ;
  RECT 1511.340 208.880 1514.880 210.000 ;
  LAYER metal1 ;
  RECT 1511.340 208.880 1514.880 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1497.700 208.880 1501.240 210.000 ;
  LAYER metal4 ;
  RECT 1497.700 208.880 1501.240 210.000 ;
  LAYER metal3 ;
  RECT 1497.700 208.880 1501.240 210.000 ;
  LAYER metal2 ;
  RECT 1497.700 208.880 1501.240 210.000 ;
  LAYER metal1 ;
  RECT 1497.700 208.880 1501.240 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1484.060 208.880 1487.600 210.000 ;
  LAYER metal4 ;
  RECT 1484.060 208.880 1487.600 210.000 ;
  LAYER metal3 ;
  RECT 1484.060 208.880 1487.600 210.000 ;
  LAYER metal2 ;
  RECT 1484.060 208.880 1487.600 210.000 ;
  LAYER metal1 ;
  RECT 1484.060 208.880 1487.600 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1417.100 208.880 1420.640 210.000 ;
  LAYER metal4 ;
  RECT 1417.100 208.880 1420.640 210.000 ;
  LAYER metal3 ;
  RECT 1417.100 208.880 1420.640 210.000 ;
  LAYER metal2 ;
  RECT 1417.100 208.880 1420.640 210.000 ;
  LAYER metal1 ;
  RECT 1417.100 208.880 1420.640 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1403.460 208.880 1407.000 210.000 ;
  LAYER metal4 ;
  RECT 1403.460 208.880 1407.000 210.000 ;
  LAYER metal3 ;
  RECT 1403.460 208.880 1407.000 210.000 ;
  LAYER metal2 ;
  RECT 1403.460 208.880 1407.000 210.000 ;
  LAYER metal1 ;
  RECT 1403.460 208.880 1407.000 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1390.440 208.880 1393.980 210.000 ;
  LAYER metal4 ;
  RECT 1390.440 208.880 1393.980 210.000 ;
  LAYER metal3 ;
  RECT 1390.440 208.880 1393.980 210.000 ;
  LAYER metal2 ;
  RECT 1390.440 208.880 1393.980 210.000 ;
  LAYER metal1 ;
  RECT 1390.440 208.880 1393.980 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1376.800 208.880 1380.340 210.000 ;
  LAYER metal4 ;
  RECT 1376.800 208.880 1380.340 210.000 ;
  LAYER metal3 ;
  RECT 1376.800 208.880 1380.340 210.000 ;
  LAYER metal2 ;
  RECT 1376.800 208.880 1380.340 210.000 ;
  LAYER metal1 ;
  RECT 1376.800 208.880 1380.340 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1363.160 208.880 1366.700 210.000 ;
  LAYER metal4 ;
  RECT 1363.160 208.880 1366.700 210.000 ;
  LAYER metal3 ;
  RECT 1363.160 208.880 1366.700 210.000 ;
  LAYER metal2 ;
  RECT 1363.160 208.880 1366.700 210.000 ;
  LAYER metal1 ;
  RECT 1363.160 208.880 1366.700 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1350.140 208.880 1353.680 210.000 ;
  LAYER metal4 ;
  RECT 1350.140 208.880 1353.680 210.000 ;
  LAYER metal3 ;
  RECT 1350.140 208.880 1353.680 210.000 ;
  LAYER metal2 ;
  RECT 1350.140 208.880 1353.680 210.000 ;
  LAYER metal1 ;
  RECT 1350.140 208.880 1353.680 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1282.560 208.880 1286.100 210.000 ;
  LAYER metal4 ;
  RECT 1282.560 208.880 1286.100 210.000 ;
  LAYER metal3 ;
  RECT 1282.560 208.880 1286.100 210.000 ;
  LAYER metal2 ;
  RECT 1282.560 208.880 1286.100 210.000 ;
  LAYER metal1 ;
  RECT 1282.560 208.880 1286.100 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1268.920 208.880 1272.460 210.000 ;
  LAYER metal4 ;
  RECT 1268.920 208.880 1272.460 210.000 ;
  LAYER metal3 ;
  RECT 1268.920 208.880 1272.460 210.000 ;
  LAYER metal2 ;
  RECT 1268.920 208.880 1272.460 210.000 ;
  LAYER metal1 ;
  RECT 1268.920 208.880 1272.460 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1255.900 208.880 1259.440 210.000 ;
  LAYER metal4 ;
  RECT 1255.900 208.880 1259.440 210.000 ;
  LAYER metal3 ;
  RECT 1255.900 208.880 1259.440 210.000 ;
  LAYER metal2 ;
  RECT 1255.900 208.880 1259.440 210.000 ;
  LAYER metal1 ;
  RECT 1255.900 208.880 1259.440 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1242.260 208.880 1245.800 210.000 ;
  LAYER metal4 ;
  RECT 1242.260 208.880 1245.800 210.000 ;
  LAYER metal3 ;
  RECT 1242.260 208.880 1245.800 210.000 ;
  LAYER metal2 ;
  RECT 1242.260 208.880 1245.800 210.000 ;
  LAYER metal1 ;
  RECT 1242.260 208.880 1245.800 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1228.620 208.880 1232.160 210.000 ;
  LAYER metal4 ;
  RECT 1228.620 208.880 1232.160 210.000 ;
  LAYER metal3 ;
  RECT 1228.620 208.880 1232.160 210.000 ;
  LAYER metal2 ;
  RECT 1228.620 208.880 1232.160 210.000 ;
  LAYER metal1 ;
  RECT 1228.620 208.880 1232.160 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1215.600 208.880 1219.140 210.000 ;
  LAYER metal4 ;
  RECT 1215.600 208.880 1219.140 210.000 ;
  LAYER metal3 ;
  RECT 1215.600 208.880 1219.140 210.000 ;
  LAYER metal2 ;
  RECT 1215.600 208.880 1219.140 210.000 ;
  LAYER metal1 ;
  RECT 1215.600 208.880 1219.140 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1148.020 208.880 1151.560 210.000 ;
  LAYER metal4 ;
  RECT 1148.020 208.880 1151.560 210.000 ;
  LAYER metal3 ;
  RECT 1148.020 208.880 1151.560 210.000 ;
  LAYER metal2 ;
  RECT 1148.020 208.880 1151.560 210.000 ;
  LAYER metal1 ;
  RECT 1148.020 208.880 1151.560 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1135.000 208.880 1138.540 210.000 ;
  LAYER metal4 ;
  RECT 1135.000 208.880 1138.540 210.000 ;
  LAYER metal3 ;
  RECT 1135.000 208.880 1138.540 210.000 ;
  LAYER metal2 ;
  RECT 1135.000 208.880 1138.540 210.000 ;
  LAYER metal1 ;
  RECT 1135.000 208.880 1138.540 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1121.360 208.880 1124.900 210.000 ;
  LAYER metal4 ;
  RECT 1121.360 208.880 1124.900 210.000 ;
  LAYER metal3 ;
  RECT 1121.360 208.880 1124.900 210.000 ;
  LAYER metal2 ;
  RECT 1121.360 208.880 1124.900 210.000 ;
  LAYER metal1 ;
  RECT 1121.360 208.880 1124.900 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1107.720 208.880 1111.260 210.000 ;
  LAYER metal4 ;
  RECT 1107.720 208.880 1111.260 210.000 ;
  LAYER metal3 ;
  RECT 1107.720 208.880 1111.260 210.000 ;
  LAYER metal2 ;
  RECT 1107.720 208.880 1111.260 210.000 ;
  LAYER metal1 ;
  RECT 1107.720 208.880 1111.260 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1094.700 208.880 1098.240 210.000 ;
  LAYER metal4 ;
  RECT 1094.700 208.880 1098.240 210.000 ;
  LAYER metal3 ;
  RECT 1094.700 208.880 1098.240 210.000 ;
  LAYER metal2 ;
  RECT 1094.700 208.880 1098.240 210.000 ;
  LAYER metal1 ;
  RECT 1094.700 208.880 1098.240 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1081.060 208.880 1084.600 210.000 ;
  LAYER metal4 ;
  RECT 1081.060 208.880 1084.600 210.000 ;
  LAYER metal3 ;
  RECT 1081.060 208.880 1084.600 210.000 ;
  LAYER metal2 ;
  RECT 1081.060 208.880 1084.600 210.000 ;
  LAYER metal1 ;
  RECT 1081.060 208.880 1084.600 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1014.100 208.880 1017.640 210.000 ;
  LAYER metal4 ;
  RECT 1014.100 208.880 1017.640 210.000 ;
  LAYER metal3 ;
  RECT 1014.100 208.880 1017.640 210.000 ;
  LAYER metal2 ;
  RECT 1014.100 208.880 1017.640 210.000 ;
  LAYER metal1 ;
  RECT 1014.100 208.880 1017.640 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1000.460 208.880 1004.000 210.000 ;
  LAYER metal4 ;
  RECT 1000.460 208.880 1004.000 210.000 ;
  LAYER metal3 ;
  RECT 1000.460 208.880 1004.000 210.000 ;
  LAYER metal2 ;
  RECT 1000.460 208.880 1004.000 210.000 ;
  LAYER metal1 ;
  RECT 1000.460 208.880 1004.000 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 986.820 208.880 990.360 210.000 ;
  LAYER metal4 ;
  RECT 986.820 208.880 990.360 210.000 ;
  LAYER metal3 ;
  RECT 986.820 208.880 990.360 210.000 ;
  LAYER metal2 ;
  RECT 986.820 208.880 990.360 210.000 ;
  LAYER metal1 ;
  RECT 986.820 208.880 990.360 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 973.800 208.880 977.340 210.000 ;
  LAYER metal4 ;
  RECT 973.800 208.880 977.340 210.000 ;
  LAYER metal3 ;
  RECT 973.800 208.880 977.340 210.000 ;
  LAYER metal2 ;
  RECT 973.800 208.880 977.340 210.000 ;
  LAYER metal1 ;
  RECT 973.800 208.880 977.340 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 960.160 208.880 963.700 210.000 ;
  LAYER metal4 ;
  RECT 960.160 208.880 963.700 210.000 ;
  LAYER metal3 ;
  RECT 960.160 208.880 963.700 210.000 ;
  LAYER metal2 ;
  RECT 960.160 208.880 963.700 210.000 ;
  LAYER metal1 ;
  RECT 960.160 208.880 963.700 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 946.520 208.880 950.060 210.000 ;
  LAYER metal4 ;
  RECT 946.520 208.880 950.060 210.000 ;
  LAYER metal3 ;
  RECT 946.520 208.880 950.060 210.000 ;
  LAYER metal2 ;
  RECT 946.520 208.880 950.060 210.000 ;
  LAYER metal1 ;
  RECT 946.520 208.880 950.060 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 879.560 208.880 883.100 210.000 ;
  LAYER metal4 ;
  RECT 879.560 208.880 883.100 210.000 ;
  LAYER metal3 ;
  RECT 879.560 208.880 883.100 210.000 ;
  LAYER metal2 ;
  RECT 879.560 208.880 883.100 210.000 ;
  LAYER metal1 ;
  RECT 879.560 208.880 883.100 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 865.920 208.880 869.460 210.000 ;
  LAYER metal4 ;
  RECT 865.920 208.880 869.460 210.000 ;
  LAYER metal3 ;
  RECT 865.920 208.880 869.460 210.000 ;
  LAYER metal2 ;
  RECT 865.920 208.880 869.460 210.000 ;
  LAYER metal1 ;
  RECT 865.920 208.880 869.460 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 852.280 208.880 855.820 210.000 ;
  LAYER metal4 ;
  RECT 852.280 208.880 855.820 210.000 ;
  LAYER metal3 ;
  RECT 852.280 208.880 855.820 210.000 ;
  LAYER metal2 ;
  RECT 852.280 208.880 855.820 210.000 ;
  LAYER metal1 ;
  RECT 852.280 208.880 855.820 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 839.260 208.880 842.800 210.000 ;
  LAYER metal4 ;
  RECT 839.260 208.880 842.800 210.000 ;
  LAYER metal3 ;
  RECT 839.260 208.880 842.800 210.000 ;
  LAYER metal2 ;
  RECT 839.260 208.880 842.800 210.000 ;
  LAYER metal1 ;
  RECT 839.260 208.880 842.800 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 825.620 208.880 829.160 210.000 ;
  LAYER metal4 ;
  RECT 825.620 208.880 829.160 210.000 ;
  LAYER metal3 ;
  RECT 825.620 208.880 829.160 210.000 ;
  LAYER metal2 ;
  RECT 825.620 208.880 829.160 210.000 ;
  LAYER metal1 ;
  RECT 825.620 208.880 829.160 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 811.980 208.880 815.520 210.000 ;
  LAYER metal4 ;
  RECT 811.980 208.880 815.520 210.000 ;
  LAYER metal3 ;
  RECT 811.980 208.880 815.520 210.000 ;
  LAYER metal2 ;
  RECT 811.980 208.880 815.520 210.000 ;
  LAYER metal1 ;
  RECT 811.980 208.880 815.520 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 745.020 208.880 748.560 210.000 ;
  LAYER metal4 ;
  RECT 745.020 208.880 748.560 210.000 ;
  LAYER metal3 ;
  RECT 745.020 208.880 748.560 210.000 ;
  LAYER metal2 ;
  RECT 745.020 208.880 748.560 210.000 ;
  LAYER metal1 ;
  RECT 745.020 208.880 748.560 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 731.380 208.880 734.920 210.000 ;
  LAYER metal4 ;
  RECT 731.380 208.880 734.920 210.000 ;
  LAYER metal3 ;
  RECT 731.380 208.880 734.920 210.000 ;
  LAYER metal2 ;
  RECT 731.380 208.880 734.920 210.000 ;
  LAYER metal1 ;
  RECT 731.380 208.880 734.920 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 718.360 208.880 721.900 210.000 ;
  LAYER metal4 ;
  RECT 718.360 208.880 721.900 210.000 ;
  LAYER metal3 ;
  RECT 718.360 208.880 721.900 210.000 ;
  LAYER metal2 ;
  RECT 718.360 208.880 721.900 210.000 ;
  LAYER metal1 ;
  RECT 718.360 208.880 721.900 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 704.720 208.880 708.260 210.000 ;
  LAYER metal4 ;
  RECT 704.720 208.880 708.260 210.000 ;
  LAYER metal3 ;
  RECT 704.720 208.880 708.260 210.000 ;
  LAYER metal2 ;
  RECT 704.720 208.880 708.260 210.000 ;
  LAYER metal1 ;
  RECT 704.720 208.880 708.260 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 691.080 208.880 694.620 210.000 ;
  LAYER metal4 ;
  RECT 691.080 208.880 694.620 210.000 ;
  LAYER metal3 ;
  RECT 691.080 208.880 694.620 210.000 ;
  LAYER metal2 ;
  RECT 691.080 208.880 694.620 210.000 ;
  LAYER metal1 ;
  RECT 691.080 208.880 694.620 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 678.060 208.880 681.600 210.000 ;
  LAYER metal4 ;
  RECT 678.060 208.880 681.600 210.000 ;
  LAYER metal3 ;
  RECT 678.060 208.880 681.600 210.000 ;
  LAYER metal2 ;
  RECT 678.060 208.880 681.600 210.000 ;
  LAYER metal1 ;
  RECT 678.060 208.880 681.600 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 610.480 208.880 614.020 210.000 ;
  LAYER metal4 ;
  RECT 610.480 208.880 614.020 210.000 ;
  LAYER metal3 ;
  RECT 610.480 208.880 614.020 210.000 ;
  LAYER metal2 ;
  RECT 610.480 208.880 614.020 210.000 ;
  LAYER metal1 ;
  RECT 610.480 208.880 614.020 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 597.460 208.880 601.000 210.000 ;
  LAYER metal4 ;
  RECT 597.460 208.880 601.000 210.000 ;
  LAYER metal3 ;
  RECT 597.460 208.880 601.000 210.000 ;
  LAYER metal2 ;
  RECT 597.460 208.880 601.000 210.000 ;
  LAYER metal1 ;
  RECT 597.460 208.880 601.000 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 583.820 208.880 587.360 210.000 ;
  LAYER metal4 ;
  RECT 583.820 208.880 587.360 210.000 ;
  LAYER metal3 ;
  RECT 583.820 208.880 587.360 210.000 ;
  LAYER metal2 ;
  RECT 583.820 208.880 587.360 210.000 ;
  LAYER metal1 ;
  RECT 583.820 208.880 587.360 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 570.180 208.880 573.720 210.000 ;
  LAYER metal4 ;
  RECT 570.180 208.880 573.720 210.000 ;
  LAYER metal3 ;
  RECT 570.180 208.880 573.720 210.000 ;
  LAYER metal2 ;
  RECT 570.180 208.880 573.720 210.000 ;
  LAYER metal1 ;
  RECT 570.180 208.880 573.720 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 557.160 208.880 560.700 210.000 ;
  LAYER metal4 ;
  RECT 557.160 208.880 560.700 210.000 ;
  LAYER metal3 ;
  RECT 557.160 208.880 560.700 210.000 ;
  LAYER metal2 ;
  RECT 557.160 208.880 560.700 210.000 ;
  LAYER metal1 ;
  RECT 557.160 208.880 560.700 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 543.520 208.880 547.060 210.000 ;
  LAYER metal4 ;
  RECT 543.520 208.880 547.060 210.000 ;
  LAYER metal3 ;
  RECT 543.520 208.880 547.060 210.000 ;
  LAYER metal2 ;
  RECT 543.520 208.880 547.060 210.000 ;
  LAYER metal1 ;
  RECT 543.520 208.880 547.060 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 475.940 208.880 479.480 210.000 ;
  LAYER metal4 ;
  RECT 475.940 208.880 479.480 210.000 ;
  LAYER metal3 ;
  RECT 475.940 208.880 479.480 210.000 ;
  LAYER metal2 ;
  RECT 475.940 208.880 479.480 210.000 ;
  LAYER metal1 ;
  RECT 475.940 208.880 479.480 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 462.920 208.880 466.460 210.000 ;
  LAYER metal4 ;
  RECT 462.920 208.880 466.460 210.000 ;
  LAYER metal3 ;
  RECT 462.920 208.880 466.460 210.000 ;
  LAYER metal2 ;
  RECT 462.920 208.880 466.460 210.000 ;
  LAYER metal1 ;
  RECT 462.920 208.880 466.460 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 449.280 208.880 452.820 210.000 ;
  LAYER metal4 ;
  RECT 449.280 208.880 452.820 210.000 ;
  LAYER metal3 ;
  RECT 449.280 208.880 452.820 210.000 ;
  LAYER metal2 ;
  RECT 449.280 208.880 452.820 210.000 ;
  LAYER metal1 ;
  RECT 449.280 208.880 452.820 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 435.640 208.880 439.180 210.000 ;
  LAYER metal4 ;
  RECT 435.640 208.880 439.180 210.000 ;
  LAYER metal3 ;
  RECT 435.640 208.880 439.180 210.000 ;
  LAYER metal2 ;
  RECT 435.640 208.880 439.180 210.000 ;
  LAYER metal1 ;
  RECT 435.640 208.880 439.180 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 422.620 208.880 426.160 210.000 ;
  LAYER metal4 ;
  RECT 422.620 208.880 426.160 210.000 ;
  LAYER metal3 ;
  RECT 422.620 208.880 426.160 210.000 ;
  LAYER metal2 ;
  RECT 422.620 208.880 426.160 210.000 ;
  LAYER metal1 ;
  RECT 422.620 208.880 426.160 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 408.980 208.880 412.520 210.000 ;
  LAYER metal4 ;
  RECT 408.980 208.880 412.520 210.000 ;
  LAYER metal3 ;
  RECT 408.980 208.880 412.520 210.000 ;
  LAYER metal2 ;
  RECT 408.980 208.880 412.520 210.000 ;
  LAYER metal1 ;
  RECT 408.980 208.880 412.520 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 342.020 208.880 345.560 210.000 ;
  LAYER metal4 ;
  RECT 342.020 208.880 345.560 210.000 ;
  LAYER metal3 ;
  RECT 342.020 208.880 345.560 210.000 ;
  LAYER metal2 ;
  RECT 342.020 208.880 345.560 210.000 ;
  LAYER metal1 ;
  RECT 342.020 208.880 345.560 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 328.380 208.880 331.920 210.000 ;
  LAYER metal4 ;
  RECT 328.380 208.880 331.920 210.000 ;
  LAYER metal3 ;
  RECT 328.380 208.880 331.920 210.000 ;
  LAYER metal2 ;
  RECT 328.380 208.880 331.920 210.000 ;
  LAYER metal1 ;
  RECT 328.380 208.880 331.920 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 314.740 208.880 318.280 210.000 ;
  LAYER metal4 ;
  RECT 314.740 208.880 318.280 210.000 ;
  LAYER metal3 ;
  RECT 314.740 208.880 318.280 210.000 ;
  LAYER metal2 ;
  RECT 314.740 208.880 318.280 210.000 ;
  LAYER metal1 ;
  RECT 314.740 208.880 318.280 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 301.720 208.880 305.260 210.000 ;
  LAYER metal4 ;
  RECT 301.720 208.880 305.260 210.000 ;
  LAYER metal3 ;
  RECT 301.720 208.880 305.260 210.000 ;
  LAYER metal2 ;
  RECT 301.720 208.880 305.260 210.000 ;
  LAYER metal1 ;
  RECT 301.720 208.880 305.260 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 288.080 208.880 291.620 210.000 ;
  LAYER metal4 ;
  RECT 288.080 208.880 291.620 210.000 ;
  LAYER metal3 ;
  RECT 288.080 208.880 291.620 210.000 ;
  LAYER metal2 ;
  RECT 288.080 208.880 291.620 210.000 ;
  LAYER metal1 ;
  RECT 288.080 208.880 291.620 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 274.440 208.880 277.980 210.000 ;
  LAYER metal4 ;
  RECT 274.440 208.880 277.980 210.000 ;
  LAYER metal3 ;
  RECT 274.440 208.880 277.980 210.000 ;
  LAYER metal2 ;
  RECT 274.440 208.880 277.980 210.000 ;
  LAYER metal1 ;
  RECT 274.440 208.880 277.980 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 207.480 208.880 211.020 210.000 ;
  LAYER metal4 ;
  RECT 207.480 208.880 211.020 210.000 ;
  LAYER metal3 ;
  RECT 207.480 208.880 211.020 210.000 ;
  LAYER metal2 ;
  RECT 207.480 208.880 211.020 210.000 ;
  LAYER metal1 ;
  RECT 207.480 208.880 211.020 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 193.840 208.880 197.380 210.000 ;
  LAYER metal4 ;
  RECT 193.840 208.880 197.380 210.000 ;
  LAYER metal3 ;
  RECT 193.840 208.880 197.380 210.000 ;
  LAYER metal2 ;
  RECT 193.840 208.880 197.380 210.000 ;
  LAYER metal1 ;
  RECT 193.840 208.880 197.380 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 180.820 208.880 184.360 210.000 ;
  LAYER metal4 ;
  RECT 180.820 208.880 184.360 210.000 ;
  LAYER metal3 ;
  RECT 180.820 208.880 184.360 210.000 ;
  LAYER metal2 ;
  RECT 180.820 208.880 184.360 210.000 ;
  LAYER metal1 ;
  RECT 180.820 208.880 184.360 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 167.180 208.880 170.720 210.000 ;
  LAYER metal4 ;
  RECT 167.180 208.880 170.720 210.000 ;
  LAYER metal3 ;
  RECT 167.180 208.880 170.720 210.000 ;
  LAYER metal2 ;
  RECT 167.180 208.880 170.720 210.000 ;
  LAYER metal1 ;
  RECT 167.180 208.880 170.720 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 153.540 208.880 157.080 210.000 ;
  LAYER metal4 ;
  RECT 153.540 208.880 157.080 210.000 ;
  LAYER metal3 ;
  RECT 153.540 208.880 157.080 210.000 ;
  LAYER metal2 ;
  RECT 153.540 208.880 157.080 210.000 ;
  LAYER metal1 ;
  RECT 153.540 208.880 157.080 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 140.520 208.880 144.060 210.000 ;
  LAYER metal4 ;
  RECT 140.520 208.880 144.060 210.000 ;
  LAYER metal3 ;
  RECT 140.520 208.880 144.060 210.000 ;
  LAYER metal2 ;
  RECT 140.520 208.880 144.060 210.000 ;
  LAYER metal1 ;
  RECT 140.520 208.880 144.060 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 72.940 208.880 76.480 210.000 ;
  LAYER metal4 ;
  RECT 72.940 208.880 76.480 210.000 ;
  LAYER metal3 ;
  RECT 72.940 208.880 76.480 210.000 ;
  LAYER metal2 ;
  RECT 72.940 208.880 76.480 210.000 ;
  LAYER metal1 ;
  RECT 72.940 208.880 76.480 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 59.300 208.880 62.840 210.000 ;
  LAYER metal4 ;
  RECT 59.300 208.880 62.840 210.000 ;
  LAYER metal3 ;
  RECT 59.300 208.880 62.840 210.000 ;
  LAYER metal2 ;
  RECT 59.300 208.880 62.840 210.000 ;
  LAYER metal1 ;
  RECT 59.300 208.880 62.840 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 46.280 208.880 49.820 210.000 ;
  LAYER metal4 ;
  RECT 46.280 208.880 49.820 210.000 ;
  LAYER metal3 ;
  RECT 46.280 208.880 49.820 210.000 ;
  LAYER metal2 ;
  RECT 46.280 208.880 49.820 210.000 ;
  LAYER metal1 ;
  RECT 46.280 208.880 49.820 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 32.640 208.880 36.180 210.000 ;
  LAYER metal4 ;
  RECT 32.640 208.880 36.180 210.000 ;
  LAYER metal3 ;
  RECT 32.640 208.880 36.180 210.000 ;
  LAYER metal2 ;
  RECT 32.640 208.880 36.180 210.000 ;
  LAYER metal1 ;
  RECT 32.640 208.880 36.180 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 19.000 208.880 22.540 210.000 ;
  LAYER metal4 ;
  RECT 19.000 208.880 22.540 210.000 ;
  LAYER metal3 ;
  RECT 19.000 208.880 22.540 210.000 ;
  LAYER metal2 ;
  RECT 19.000 208.880 22.540 210.000 ;
  LAYER metal1 ;
  RECT 19.000 208.880 22.540 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 7.220 208.880 10.760 210.000 ;
  LAYER metal4 ;
  RECT 7.220 208.880 10.760 210.000 ;
  LAYER metal3 ;
  RECT 7.220 208.880 10.760 210.000 ;
  LAYER metal2 ;
  RECT 7.220 208.880 10.760 210.000 ;
  LAYER metal1 ;
  RECT 7.220 208.880 10.760 210.000 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3559.820 0.000 3563.360 1.120 ;
  LAYER metal4 ;
  RECT 3559.820 0.000 3563.360 1.120 ;
  LAYER metal3 ;
  RECT 3559.820 0.000 3563.360 1.120 ;
  LAYER metal2 ;
  RECT 3559.820 0.000 3563.360 1.120 ;
  LAYER metal1 ;
  RECT 3559.820 0.000 3563.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3551.140 0.000 3554.680 1.120 ;
  LAYER metal4 ;
  RECT 3551.140 0.000 3554.680 1.120 ;
  LAYER metal3 ;
  RECT 3551.140 0.000 3554.680 1.120 ;
  LAYER metal2 ;
  RECT 3551.140 0.000 3554.680 1.120 ;
  LAYER metal1 ;
  RECT 3551.140 0.000 3554.680 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3537.500 0.000 3541.040 1.120 ;
  LAYER metal4 ;
  RECT 3537.500 0.000 3541.040 1.120 ;
  LAYER metal3 ;
  RECT 3537.500 0.000 3541.040 1.120 ;
  LAYER metal2 ;
  RECT 3537.500 0.000 3541.040 1.120 ;
  LAYER metal1 ;
  RECT 3537.500 0.000 3541.040 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3524.480 0.000 3528.020 1.120 ;
  LAYER metal4 ;
  RECT 3524.480 0.000 3528.020 1.120 ;
  LAYER metal3 ;
  RECT 3524.480 0.000 3528.020 1.120 ;
  LAYER metal2 ;
  RECT 3524.480 0.000 3528.020 1.120 ;
  LAYER metal1 ;
  RECT 3524.480 0.000 3528.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3456.900 0.000 3460.440 1.120 ;
  LAYER metal4 ;
  RECT 3456.900 0.000 3460.440 1.120 ;
  LAYER metal3 ;
  RECT 3456.900 0.000 3460.440 1.120 ;
  LAYER metal2 ;
  RECT 3456.900 0.000 3460.440 1.120 ;
  LAYER metal1 ;
  RECT 3456.900 0.000 3460.440 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3443.260 0.000 3446.800 1.120 ;
  LAYER metal4 ;
  RECT 3443.260 0.000 3446.800 1.120 ;
  LAYER metal3 ;
  RECT 3443.260 0.000 3446.800 1.120 ;
  LAYER metal2 ;
  RECT 3443.260 0.000 3446.800 1.120 ;
  LAYER metal1 ;
  RECT 3443.260 0.000 3446.800 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3430.240 0.000 3433.780 1.120 ;
  LAYER metal4 ;
  RECT 3430.240 0.000 3433.780 1.120 ;
  LAYER metal3 ;
  RECT 3430.240 0.000 3433.780 1.120 ;
  LAYER metal2 ;
  RECT 3430.240 0.000 3433.780 1.120 ;
  LAYER metal1 ;
  RECT 3430.240 0.000 3433.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3416.600 0.000 3420.140 1.120 ;
  LAYER metal4 ;
  RECT 3416.600 0.000 3420.140 1.120 ;
  LAYER metal3 ;
  RECT 3416.600 0.000 3420.140 1.120 ;
  LAYER metal2 ;
  RECT 3416.600 0.000 3420.140 1.120 ;
  LAYER metal1 ;
  RECT 3416.600 0.000 3420.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3402.960 0.000 3406.500 1.120 ;
  LAYER metal4 ;
  RECT 3402.960 0.000 3406.500 1.120 ;
  LAYER metal3 ;
  RECT 3402.960 0.000 3406.500 1.120 ;
  LAYER metal2 ;
  RECT 3402.960 0.000 3406.500 1.120 ;
  LAYER metal1 ;
  RECT 3402.960 0.000 3406.500 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3389.940 0.000 3393.480 1.120 ;
  LAYER metal4 ;
  RECT 3389.940 0.000 3393.480 1.120 ;
  LAYER metal3 ;
  RECT 3389.940 0.000 3393.480 1.120 ;
  LAYER metal2 ;
  RECT 3389.940 0.000 3393.480 1.120 ;
  LAYER metal1 ;
  RECT 3389.940 0.000 3393.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3322.360 0.000 3325.900 1.120 ;
  LAYER metal4 ;
  RECT 3322.360 0.000 3325.900 1.120 ;
  LAYER metal3 ;
  RECT 3322.360 0.000 3325.900 1.120 ;
  LAYER metal2 ;
  RECT 3322.360 0.000 3325.900 1.120 ;
  LAYER metal1 ;
  RECT 3322.360 0.000 3325.900 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3309.340 0.000 3312.880 1.120 ;
  LAYER metal4 ;
  RECT 3309.340 0.000 3312.880 1.120 ;
  LAYER metal3 ;
  RECT 3309.340 0.000 3312.880 1.120 ;
  LAYER metal2 ;
  RECT 3309.340 0.000 3312.880 1.120 ;
  LAYER metal1 ;
  RECT 3309.340 0.000 3312.880 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3295.700 0.000 3299.240 1.120 ;
  LAYER metal4 ;
  RECT 3295.700 0.000 3299.240 1.120 ;
  LAYER metal3 ;
  RECT 3295.700 0.000 3299.240 1.120 ;
  LAYER metal2 ;
  RECT 3295.700 0.000 3299.240 1.120 ;
  LAYER metal1 ;
  RECT 3295.700 0.000 3299.240 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3282.060 0.000 3285.600 1.120 ;
  LAYER metal4 ;
  RECT 3282.060 0.000 3285.600 1.120 ;
  LAYER metal3 ;
  RECT 3282.060 0.000 3285.600 1.120 ;
  LAYER metal2 ;
  RECT 3282.060 0.000 3285.600 1.120 ;
  LAYER metal1 ;
  RECT 3282.060 0.000 3285.600 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3269.040 0.000 3272.580 1.120 ;
  LAYER metal4 ;
  RECT 3269.040 0.000 3272.580 1.120 ;
  LAYER metal3 ;
  RECT 3269.040 0.000 3272.580 1.120 ;
  LAYER metal2 ;
  RECT 3269.040 0.000 3272.580 1.120 ;
  LAYER metal1 ;
  RECT 3269.040 0.000 3272.580 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3255.400 0.000 3258.940 1.120 ;
  LAYER metal4 ;
  RECT 3255.400 0.000 3258.940 1.120 ;
  LAYER metal3 ;
  RECT 3255.400 0.000 3258.940 1.120 ;
  LAYER metal2 ;
  RECT 3255.400 0.000 3258.940 1.120 ;
  LAYER metal1 ;
  RECT 3255.400 0.000 3258.940 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3188.440 0.000 3191.980 1.120 ;
  LAYER metal4 ;
  RECT 3188.440 0.000 3191.980 1.120 ;
  LAYER metal3 ;
  RECT 3188.440 0.000 3191.980 1.120 ;
  LAYER metal2 ;
  RECT 3188.440 0.000 3191.980 1.120 ;
  LAYER metal1 ;
  RECT 3188.440 0.000 3191.980 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3174.800 0.000 3178.340 1.120 ;
  LAYER metal4 ;
  RECT 3174.800 0.000 3178.340 1.120 ;
  LAYER metal3 ;
  RECT 3174.800 0.000 3178.340 1.120 ;
  LAYER metal2 ;
  RECT 3174.800 0.000 3178.340 1.120 ;
  LAYER metal1 ;
  RECT 3174.800 0.000 3178.340 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3161.160 0.000 3164.700 1.120 ;
  LAYER metal4 ;
  RECT 3161.160 0.000 3164.700 1.120 ;
  LAYER metal3 ;
  RECT 3161.160 0.000 3164.700 1.120 ;
  LAYER metal2 ;
  RECT 3161.160 0.000 3164.700 1.120 ;
  LAYER metal1 ;
  RECT 3161.160 0.000 3164.700 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3148.140 0.000 3151.680 1.120 ;
  LAYER metal4 ;
  RECT 3148.140 0.000 3151.680 1.120 ;
  LAYER metal3 ;
  RECT 3148.140 0.000 3151.680 1.120 ;
  LAYER metal2 ;
  RECT 3148.140 0.000 3151.680 1.120 ;
  LAYER metal1 ;
  RECT 3148.140 0.000 3151.680 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3134.500 0.000 3138.040 1.120 ;
  LAYER metal4 ;
  RECT 3134.500 0.000 3138.040 1.120 ;
  LAYER metal3 ;
  RECT 3134.500 0.000 3138.040 1.120 ;
  LAYER metal2 ;
  RECT 3134.500 0.000 3138.040 1.120 ;
  LAYER metal1 ;
  RECT 3134.500 0.000 3138.040 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3120.860 0.000 3124.400 1.120 ;
  LAYER metal4 ;
  RECT 3120.860 0.000 3124.400 1.120 ;
  LAYER metal3 ;
  RECT 3120.860 0.000 3124.400 1.120 ;
  LAYER metal2 ;
  RECT 3120.860 0.000 3124.400 1.120 ;
  LAYER metal1 ;
  RECT 3120.860 0.000 3124.400 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3053.900 0.000 3057.440 1.120 ;
  LAYER metal4 ;
  RECT 3053.900 0.000 3057.440 1.120 ;
  LAYER metal3 ;
  RECT 3053.900 0.000 3057.440 1.120 ;
  LAYER metal2 ;
  RECT 3053.900 0.000 3057.440 1.120 ;
  LAYER metal1 ;
  RECT 3053.900 0.000 3057.440 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3040.260 0.000 3043.800 1.120 ;
  LAYER metal4 ;
  RECT 3040.260 0.000 3043.800 1.120 ;
  LAYER metal3 ;
  RECT 3040.260 0.000 3043.800 1.120 ;
  LAYER metal2 ;
  RECT 3040.260 0.000 3043.800 1.120 ;
  LAYER metal1 ;
  RECT 3040.260 0.000 3043.800 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3026.620 0.000 3030.160 1.120 ;
  LAYER metal4 ;
  RECT 3026.620 0.000 3030.160 1.120 ;
  LAYER metal3 ;
  RECT 3026.620 0.000 3030.160 1.120 ;
  LAYER metal2 ;
  RECT 3026.620 0.000 3030.160 1.120 ;
  LAYER metal1 ;
  RECT 3026.620 0.000 3030.160 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 3013.600 0.000 3017.140 1.120 ;
  LAYER metal4 ;
  RECT 3013.600 0.000 3017.140 1.120 ;
  LAYER metal3 ;
  RECT 3013.600 0.000 3017.140 1.120 ;
  LAYER metal2 ;
  RECT 3013.600 0.000 3017.140 1.120 ;
  LAYER metal1 ;
  RECT 3013.600 0.000 3017.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2999.960 0.000 3003.500 1.120 ;
  LAYER metal4 ;
  RECT 2999.960 0.000 3003.500 1.120 ;
  LAYER metal3 ;
  RECT 2999.960 0.000 3003.500 1.120 ;
  LAYER metal2 ;
  RECT 2999.960 0.000 3003.500 1.120 ;
  LAYER metal1 ;
  RECT 2999.960 0.000 3003.500 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2986.320 0.000 2989.860 1.120 ;
  LAYER metal4 ;
  RECT 2986.320 0.000 2989.860 1.120 ;
  LAYER metal3 ;
  RECT 2986.320 0.000 2989.860 1.120 ;
  LAYER metal2 ;
  RECT 2986.320 0.000 2989.860 1.120 ;
  LAYER metal1 ;
  RECT 2986.320 0.000 2989.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2919.360 0.000 2922.900 1.120 ;
  LAYER metal4 ;
  RECT 2919.360 0.000 2922.900 1.120 ;
  LAYER metal3 ;
  RECT 2919.360 0.000 2922.900 1.120 ;
  LAYER metal2 ;
  RECT 2919.360 0.000 2922.900 1.120 ;
  LAYER metal1 ;
  RECT 2919.360 0.000 2922.900 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2905.720 0.000 2909.260 1.120 ;
  LAYER metal4 ;
  RECT 2905.720 0.000 2909.260 1.120 ;
  LAYER metal3 ;
  RECT 2905.720 0.000 2909.260 1.120 ;
  LAYER metal2 ;
  RECT 2905.720 0.000 2909.260 1.120 ;
  LAYER metal1 ;
  RECT 2905.720 0.000 2909.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2892.700 0.000 2896.240 1.120 ;
  LAYER metal4 ;
  RECT 2892.700 0.000 2896.240 1.120 ;
  LAYER metal3 ;
  RECT 2892.700 0.000 2896.240 1.120 ;
  LAYER metal2 ;
  RECT 2892.700 0.000 2896.240 1.120 ;
  LAYER metal1 ;
  RECT 2892.700 0.000 2896.240 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2879.060 0.000 2882.600 1.120 ;
  LAYER metal4 ;
  RECT 2879.060 0.000 2882.600 1.120 ;
  LAYER metal3 ;
  RECT 2879.060 0.000 2882.600 1.120 ;
  LAYER metal2 ;
  RECT 2879.060 0.000 2882.600 1.120 ;
  LAYER metal1 ;
  RECT 2879.060 0.000 2882.600 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2865.420 0.000 2868.960 1.120 ;
  LAYER metal4 ;
  RECT 2865.420 0.000 2868.960 1.120 ;
  LAYER metal3 ;
  RECT 2865.420 0.000 2868.960 1.120 ;
  LAYER metal2 ;
  RECT 2865.420 0.000 2868.960 1.120 ;
  LAYER metal1 ;
  RECT 2865.420 0.000 2868.960 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2852.400 0.000 2855.940 1.120 ;
  LAYER metal4 ;
  RECT 2852.400 0.000 2855.940 1.120 ;
  LAYER metal3 ;
  RECT 2852.400 0.000 2855.940 1.120 ;
  LAYER metal2 ;
  RECT 2852.400 0.000 2855.940 1.120 ;
  LAYER metal1 ;
  RECT 2852.400 0.000 2855.940 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2784.820 0.000 2788.360 1.120 ;
  LAYER metal4 ;
  RECT 2784.820 0.000 2788.360 1.120 ;
  LAYER metal3 ;
  RECT 2784.820 0.000 2788.360 1.120 ;
  LAYER metal2 ;
  RECT 2784.820 0.000 2788.360 1.120 ;
  LAYER metal1 ;
  RECT 2784.820 0.000 2788.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2771.800 0.000 2775.340 1.120 ;
  LAYER metal4 ;
  RECT 2771.800 0.000 2775.340 1.120 ;
  LAYER metal3 ;
  RECT 2771.800 0.000 2775.340 1.120 ;
  LAYER metal2 ;
  RECT 2771.800 0.000 2775.340 1.120 ;
  LAYER metal1 ;
  RECT 2771.800 0.000 2775.340 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2758.160 0.000 2761.700 1.120 ;
  LAYER metal4 ;
  RECT 2758.160 0.000 2761.700 1.120 ;
  LAYER metal3 ;
  RECT 2758.160 0.000 2761.700 1.120 ;
  LAYER metal2 ;
  RECT 2758.160 0.000 2761.700 1.120 ;
  LAYER metal1 ;
  RECT 2758.160 0.000 2761.700 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2744.520 0.000 2748.060 1.120 ;
  LAYER metal4 ;
  RECT 2744.520 0.000 2748.060 1.120 ;
  LAYER metal3 ;
  RECT 2744.520 0.000 2748.060 1.120 ;
  LAYER metal2 ;
  RECT 2744.520 0.000 2748.060 1.120 ;
  LAYER metal1 ;
  RECT 2744.520 0.000 2748.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2731.500 0.000 2735.040 1.120 ;
  LAYER metal4 ;
  RECT 2731.500 0.000 2735.040 1.120 ;
  LAYER metal3 ;
  RECT 2731.500 0.000 2735.040 1.120 ;
  LAYER metal2 ;
  RECT 2731.500 0.000 2735.040 1.120 ;
  LAYER metal1 ;
  RECT 2731.500 0.000 2735.040 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2717.860 0.000 2721.400 1.120 ;
  LAYER metal4 ;
  RECT 2717.860 0.000 2721.400 1.120 ;
  LAYER metal3 ;
  RECT 2717.860 0.000 2721.400 1.120 ;
  LAYER metal2 ;
  RECT 2717.860 0.000 2721.400 1.120 ;
  LAYER metal1 ;
  RECT 2717.860 0.000 2721.400 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2650.900 0.000 2654.440 1.120 ;
  LAYER metal4 ;
  RECT 2650.900 0.000 2654.440 1.120 ;
  LAYER metal3 ;
  RECT 2650.900 0.000 2654.440 1.120 ;
  LAYER metal2 ;
  RECT 2650.900 0.000 2654.440 1.120 ;
  LAYER metal1 ;
  RECT 2650.900 0.000 2654.440 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2637.260 0.000 2640.800 1.120 ;
  LAYER metal4 ;
  RECT 2637.260 0.000 2640.800 1.120 ;
  LAYER metal3 ;
  RECT 2637.260 0.000 2640.800 1.120 ;
  LAYER metal2 ;
  RECT 2637.260 0.000 2640.800 1.120 ;
  LAYER metal1 ;
  RECT 2637.260 0.000 2640.800 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2623.620 0.000 2627.160 1.120 ;
  LAYER metal4 ;
  RECT 2623.620 0.000 2627.160 1.120 ;
  LAYER metal3 ;
  RECT 2623.620 0.000 2627.160 1.120 ;
  LAYER metal2 ;
  RECT 2623.620 0.000 2627.160 1.120 ;
  LAYER metal1 ;
  RECT 2623.620 0.000 2627.160 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2609.980 0.000 2613.520 1.120 ;
  LAYER metal4 ;
  RECT 2609.980 0.000 2613.520 1.120 ;
  LAYER metal3 ;
  RECT 2609.980 0.000 2613.520 1.120 ;
  LAYER metal2 ;
  RECT 2609.980 0.000 2613.520 1.120 ;
  LAYER metal1 ;
  RECT 2609.980 0.000 2613.520 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2596.960 0.000 2600.500 1.120 ;
  LAYER metal4 ;
  RECT 2596.960 0.000 2600.500 1.120 ;
  LAYER metal3 ;
  RECT 2596.960 0.000 2600.500 1.120 ;
  LAYER metal2 ;
  RECT 2596.960 0.000 2600.500 1.120 ;
  LAYER metal1 ;
  RECT 2596.960 0.000 2600.500 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2583.320 0.000 2586.860 1.120 ;
  LAYER metal4 ;
  RECT 2583.320 0.000 2586.860 1.120 ;
  LAYER metal3 ;
  RECT 2583.320 0.000 2586.860 1.120 ;
  LAYER metal2 ;
  RECT 2583.320 0.000 2586.860 1.120 ;
  LAYER metal1 ;
  RECT 2583.320 0.000 2586.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2516.360 0.000 2519.900 1.120 ;
  LAYER metal4 ;
  RECT 2516.360 0.000 2519.900 1.120 ;
  LAYER metal3 ;
  RECT 2516.360 0.000 2519.900 1.120 ;
  LAYER metal2 ;
  RECT 2516.360 0.000 2519.900 1.120 ;
  LAYER metal1 ;
  RECT 2516.360 0.000 2519.900 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2502.720 0.000 2506.260 1.120 ;
  LAYER metal4 ;
  RECT 2502.720 0.000 2506.260 1.120 ;
  LAYER metal3 ;
  RECT 2502.720 0.000 2506.260 1.120 ;
  LAYER metal2 ;
  RECT 2502.720 0.000 2506.260 1.120 ;
  LAYER metal1 ;
  RECT 2502.720 0.000 2506.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2489.080 0.000 2492.620 1.120 ;
  LAYER metal4 ;
  RECT 2489.080 0.000 2492.620 1.120 ;
  LAYER metal3 ;
  RECT 2489.080 0.000 2492.620 1.120 ;
  LAYER metal2 ;
  RECT 2489.080 0.000 2492.620 1.120 ;
  LAYER metal1 ;
  RECT 2489.080 0.000 2492.620 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2476.060 0.000 2479.600 1.120 ;
  LAYER metal4 ;
  RECT 2476.060 0.000 2479.600 1.120 ;
  LAYER metal3 ;
  RECT 2476.060 0.000 2479.600 1.120 ;
  LAYER metal2 ;
  RECT 2476.060 0.000 2479.600 1.120 ;
  LAYER metal1 ;
  RECT 2476.060 0.000 2479.600 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2462.420 0.000 2465.960 1.120 ;
  LAYER metal4 ;
  RECT 2462.420 0.000 2465.960 1.120 ;
  LAYER metal3 ;
  RECT 2462.420 0.000 2465.960 1.120 ;
  LAYER metal2 ;
  RECT 2462.420 0.000 2465.960 1.120 ;
  LAYER metal1 ;
  RECT 2462.420 0.000 2465.960 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2448.780 0.000 2452.320 1.120 ;
  LAYER metal4 ;
  RECT 2448.780 0.000 2452.320 1.120 ;
  LAYER metal3 ;
  RECT 2448.780 0.000 2452.320 1.120 ;
  LAYER metal2 ;
  RECT 2448.780 0.000 2452.320 1.120 ;
  LAYER metal1 ;
  RECT 2448.780 0.000 2452.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2381.820 0.000 2385.360 1.120 ;
  LAYER metal4 ;
  RECT 2381.820 0.000 2385.360 1.120 ;
  LAYER metal3 ;
  RECT 2381.820 0.000 2385.360 1.120 ;
  LAYER metal2 ;
  RECT 2381.820 0.000 2385.360 1.120 ;
  LAYER metal1 ;
  RECT 2381.820 0.000 2385.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2368.180 0.000 2371.720 1.120 ;
  LAYER metal4 ;
  RECT 2368.180 0.000 2371.720 1.120 ;
  LAYER metal3 ;
  RECT 2368.180 0.000 2371.720 1.120 ;
  LAYER metal2 ;
  RECT 2368.180 0.000 2371.720 1.120 ;
  LAYER metal1 ;
  RECT 2368.180 0.000 2371.720 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2355.160 0.000 2358.700 1.120 ;
  LAYER metal4 ;
  RECT 2355.160 0.000 2358.700 1.120 ;
  LAYER metal3 ;
  RECT 2355.160 0.000 2358.700 1.120 ;
  LAYER metal2 ;
  RECT 2355.160 0.000 2358.700 1.120 ;
  LAYER metal1 ;
  RECT 2355.160 0.000 2358.700 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2341.520 0.000 2345.060 1.120 ;
  LAYER metal4 ;
  RECT 2341.520 0.000 2345.060 1.120 ;
  LAYER metal3 ;
  RECT 2341.520 0.000 2345.060 1.120 ;
  LAYER metal2 ;
  RECT 2341.520 0.000 2345.060 1.120 ;
  LAYER metal1 ;
  RECT 2341.520 0.000 2345.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2327.880 0.000 2331.420 1.120 ;
  LAYER metal4 ;
  RECT 2327.880 0.000 2331.420 1.120 ;
  LAYER metal3 ;
  RECT 2327.880 0.000 2331.420 1.120 ;
  LAYER metal2 ;
  RECT 2327.880 0.000 2331.420 1.120 ;
  LAYER metal1 ;
  RECT 2327.880 0.000 2331.420 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2314.860 0.000 2318.400 1.120 ;
  LAYER metal4 ;
  RECT 2314.860 0.000 2318.400 1.120 ;
  LAYER metal3 ;
  RECT 2314.860 0.000 2318.400 1.120 ;
  LAYER metal2 ;
  RECT 2314.860 0.000 2318.400 1.120 ;
  LAYER metal1 ;
  RECT 2314.860 0.000 2318.400 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2247.280 0.000 2250.820 1.120 ;
  LAYER metal4 ;
  RECT 2247.280 0.000 2250.820 1.120 ;
  LAYER metal3 ;
  RECT 2247.280 0.000 2250.820 1.120 ;
  LAYER metal2 ;
  RECT 2247.280 0.000 2250.820 1.120 ;
  LAYER metal1 ;
  RECT 2247.280 0.000 2250.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2234.260 0.000 2237.800 1.120 ;
  LAYER metal4 ;
  RECT 2234.260 0.000 2237.800 1.120 ;
  LAYER metal3 ;
  RECT 2234.260 0.000 2237.800 1.120 ;
  LAYER metal2 ;
  RECT 2234.260 0.000 2237.800 1.120 ;
  LAYER metal1 ;
  RECT 2234.260 0.000 2237.800 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2220.620 0.000 2224.160 1.120 ;
  LAYER metal4 ;
  RECT 2220.620 0.000 2224.160 1.120 ;
  LAYER metal3 ;
  RECT 2220.620 0.000 2224.160 1.120 ;
  LAYER metal2 ;
  RECT 2220.620 0.000 2224.160 1.120 ;
  LAYER metal1 ;
  RECT 2220.620 0.000 2224.160 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2206.980 0.000 2210.520 1.120 ;
  LAYER metal4 ;
  RECT 2206.980 0.000 2210.520 1.120 ;
  LAYER metal3 ;
  RECT 2206.980 0.000 2210.520 1.120 ;
  LAYER metal2 ;
  RECT 2206.980 0.000 2210.520 1.120 ;
  LAYER metal1 ;
  RECT 2206.980 0.000 2210.520 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2193.340 0.000 2196.880 1.120 ;
  LAYER metal4 ;
  RECT 2193.340 0.000 2196.880 1.120 ;
  LAYER metal3 ;
  RECT 2193.340 0.000 2196.880 1.120 ;
  LAYER metal2 ;
  RECT 2193.340 0.000 2196.880 1.120 ;
  LAYER metal1 ;
  RECT 2193.340 0.000 2196.880 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2180.320 0.000 2183.860 1.120 ;
  LAYER metal4 ;
  RECT 2180.320 0.000 2183.860 1.120 ;
  LAYER metal3 ;
  RECT 2180.320 0.000 2183.860 1.120 ;
  LAYER metal2 ;
  RECT 2180.320 0.000 2183.860 1.120 ;
  LAYER metal1 ;
  RECT 2180.320 0.000 2183.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2112.740 0.000 2116.280 1.120 ;
  LAYER metal4 ;
  RECT 2112.740 0.000 2116.280 1.120 ;
  LAYER metal3 ;
  RECT 2112.740 0.000 2116.280 1.120 ;
  LAYER metal2 ;
  RECT 2112.740 0.000 2116.280 1.120 ;
  LAYER metal1 ;
  RECT 2112.740 0.000 2116.280 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2099.720 0.000 2103.260 1.120 ;
  LAYER metal4 ;
  RECT 2099.720 0.000 2103.260 1.120 ;
  LAYER metal3 ;
  RECT 2099.720 0.000 2103.260 1.120 ;
  LAYER metal2 ;
  RECT 2099.720 0.000 2103.260 1.120 ;
  LAYER metal1 ;
  RECT 2099.720 0.000 2103.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2086.080 0.000 2089.620 1.120 ;
  LAYER metal4 ;
  RECT 2086.080 0.000 2089.620 1.120 ;
  LAYER metal3 ;
  RECT 2086.080 0.000 2089.620 1.120 ;
  LAYER metal2 ;
  RECT 2086.080 0.000 2089.620 1.120 ;
  LAYER metal1 ;
  RECT 2086.080 0.000 2089.620 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2072.440 0.000 2075.980 1.120 ;
  LAYER metal4 ;
  RECT 2072.440 0.000 2075.980 1.120 ;
  LAYER metal3 ;
  RECT 2072.440 0.000 2075.980 1.120 ;
  LAYER metal2 ;
  RECT 2072.440 0.000 2075.980 1.120 ;
  LAYER metal1 ;
  RECT 2072.440 0.000 2075.980 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2059.420 0.000 2062.960 1.120 ;
  LAYER metal4 ;
  RECT 2059.420 0.000 2062.960 1.120 ;
  LAYER metal3 ;
  RECT 2059.420 0.000 2062.960 1.120 ;
  LAYER metal2 ;
  RECT 2059.420 0.000 2062.960 1.120 ;
  LAYER metal1 ;
  RECT 2059.420 0.000 2062.960 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 2045.780 0.000 2049.320 1.120 ;
  LAYER metal4 ;
  RECT 2045.780 0.000 2049.320 1.120 ;
  LAYER metal3 ;
  RECT 2045.780 0.000 2049.320 1.120 ;
  LAYER metal2 ;
  RECT 2045.780 0.000 2049.320 1.120 ;
  LAYER metal1 ;
  RECT 2045.780 0.000 2049.320 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1978.820 0.000 1982.360 1.120 ;
  LAYER metal4 ;
  RECT 1978.820 0.000 1982.360 1.120 ;
  LAYER metal3 ;
  RECT 1978.820 0.000 1982.360 1.120 ;
  LAYER metal2 ;
  RECT 1978.820 0.000 1982.360 1.120 ;
  LAYER metal1 ;
  RECT 1978.820 0.000 1982.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1965.180 0.000 1968.720 1.120 ;
  LAYER metal4 ;
  RECT 1965.180 0.000 1968.720 1.120 ;
  LAYER metal3 ;
  RECT 1965.180 0.000 1968.720 1.120 ;
  LAYER metal2 ;
  RECT 1965.180 0.000 1968.720 1.120 ;
  LAYER metal1 ;
  RECT 1965.180 0.000 1968.720 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1951.540 0.000 1955.080 1.120 ;
  LAYER metal4 ;
  RECT 1951.540 0.000 1955.080 1.120 ;
  LAYER metal3 ;
  RECT 1951.540 0.000 1955.080 1.120 ;
  LAYER metal2 ;
  RECT 1951.540 0.000 1955.080 1.120 ;
  LAYER metal1 ;
  RECT 1951.540 0.000 1955.080 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1938.520 0.000 1942.060 1.120 ;
  LAYER metal4 ;
  RECT 1938.520 0.000 1942.060 1.120 ;
  LAYER metal3 ;
  RECT 1938.520 0.000 1942.060 1.120 ;
  LAYER metal2 ;
  RECT 1938.520 0.000 1942.060 1.120 ;
  LAYER metal1 ;
  RECT 1938.520 0.000 1942.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1924.880 0.000 1928.420 1.120 ;
  LAYER metal4 ;
  RECT 1924.880 0.000 1928.420 1.120 ;
  LAYER metal3 ;
  RECT 1924.880 0.000 1928.420 1.120 ;
  LAYER metal2 ;
  RECT 1924.880 0.000 1928.420 1.120 ;
  LAYER metal1 ;
  RECT 1924.880 0.000 1928.420 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1911.240 0.000 1914.780 1.120 ;
  LAYER metal4 ;
  RECT 1911.240 0.000 1914.780 1.120 ;
  LAYER metal3 ;
  RECT 1911.240 0.000 1914.780 1.120 ;
  LAYER metal2 ;
  RECT 1911.240 0.000 1914.780 1.120 ;
  LAYER metal1 ;
  RECT 1911.240 0.000 1914.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1844.280 0.000 1847.820 1.120 ;
  LAYER metal4 ;
  RECT 1844.280 0.000 1847.820 1.120 ;
  LAYER metal3 ;
  RECT 1844.280 0.000 1847.820 1.120 ;
  LAYER metal2 ;
  RECT 1844.280 0.000 1847.820 1.120 ;
  LAYER metal1 ;
  RECT 1844.280 0.000 1847.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1830.640 0.000 1834.180 1.120 ;
  LAYER metal4 ;
  RECT 1830.640 0.000 1834.180 1.120 ;
  LAYER metal3 ;
  RECT 1830.640 0.000 1834.180 1.120 ;
  LAYER metal2 ;
  RECT 1830.640 0.000 1834.180 1.120 ;
  LAYER metal1 ;
  RECT 1830.640 0.000 1834.180 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1821.960 0.000 1825.500 1.120 ;
  LAYER metal4 ;
  RECT 1821.960 0.000 1825.500 1.120 ;
  LAYER metal3 ;
  RECT 1821.960 0.000 1825.500 1.120 ;
  LAYER metal2 ;
  RECT 1821.960 0.000 1825.500 1.120 ;
  LAYER metal1 ;
  RECT 1821.960 0.000 1825.500 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1808.320 0.000 1811.860 1.120 ;
  LAYER metal4 ;
  RECT 1808.320 0.000 1811.860 1.120 ;
  LAYER metal3 ;
  RECT 1808.320 0.000 1811.860 1.120 ;
  LAYER metal2 ;
  RECT 1808.320 0.000 1811.860 1.120 ;
  LAYER metal1 ;
  RECT 1808.320 0.000 1811.860 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1779.800 0.000 1783.340 1.120 ;
  LAYER metal4 ;
  RECT 1779.800 0.000 1783.340 1.120 ;
  LAYER metal3 ;
  RECT 1779.800 0.000 1783.340 1.120 ;
  LAYER metal2 ;
  RECT 1779.800 0.000 1783.340 1.120 ;
  LAYER metal1 ;
  RECT 1779.800 0.000 1783.340 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1754.380 0.000 1757.920 1.120 ;
  LAYER metal4 ;
  RECT 1754.380 0.000 1757.920 1.120 ;
  LAYER metal3 ;
  RECT 1754.380 0.000 1757.920 1.120 ;
  LAYER metal2 ;
  RECT 1754.380 0.000 1757.920 1.120 ;
  LAYER metal1 ;
  RECT 1754.380 0.000 1757.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1685.560 0.000 1689.100 1.120 ;
  LAYER metal4 ;
  RECT 1685.560 0.000 1689.100 1.120 ;
  LAYER metal3 ;
  RECT 1685.560 0.000 1689.100 1.120 ;
  LAYER metal2 ;
  RECT 1685.560 0.000 1689.100 1.120 ;
  LAYER metal1 ;
  RECT 1685.560 0.000 1689.100 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1672.540 0.000 1676.080 1.120 ;
  LAYER metal4 ;
  RECT 1672.540 0.000 1676.080 1.120 ;
  LAYER metal3 ;
  RECT 1672.540 0.000 1676.080 1.120 ;
  LAYER metal2 ;
  RECT 1672.540 0.000 1676.080 1.120 ;
  LAYER metal1 ;
  RECT 1672.540 0.000 1676.080 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1658.900 0.000 1662.440 1.120 ;
  LAYER metal4 ;
  RECT 1658.900 0.000 1662.440 1.120 ;
  LAYER metal3 ;
  RECT 1658.900 0.000 1662.440 1.120 ;
  LAYER metal2 ;
  RECT 1658.900 0.000 1662.440 1.120 ;
  LAYER metal1 ;
  RECT 1658.900 0.000 1662.440 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1645.260 0.000 1648.800 1.120 ;
  LAYER metal4 ;
  RECT 1645.260 0.000 1648.800 1.120 ;
  LAYER metal3 ;
  RECT 1645.260 0.000 1648.800 1.120 ;
  LAYER metal2 ;
  RECT 1645.260 0.000 1648.800 1.120 ;
  LAYER metal1 ;
  RECT 1645.260 0.000 1648.800 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1632.240 0.000 1635.780 1.120 ;
  LAYER metal4 ;
  RECT 1632.240 0.000 1635.780 1.120 ;
  LAYER metal3 ;
  RECT 1632.240 0.000 1635.780 1.120 ;
  LAYER metal2 ;
  RECT 1632.240 0.000 1635.780 1.120 ;
  LAYER metal1 ;
  RECT 1632.240 0.000 1635.780 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1618.600 0.000 1622.140 1.120 ;
  LAYER metal4 ;
  RECT 1618.600 0.000 1622.140 1.120 ;
  LAYER metal3 ;
  RECT 1618.600 0.000 1622.140 1.120 ;
  LAYER metal2 ;
  RECT 1618.600 0.000 1622.140 1.120 ;
  LAYER metal1 ;
  RECT 1618.600 0.000 1622.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1551.640 0.000 1555.180 1.120 ;
  LAYER metal4 ;
  RECT 1551.640 0.000 1555.180 1.120 ;
  LAYER metal3 ;
  RECT 1551.640 0.000 1555.180 1.120 ;
  LAYER metal2 ;
  RECT 1551.640 0.000 1555.180 1.120 ;
  LAYER metal1 ;
  RECT 1551.640 0.000 1555.180 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1538.000 0.000 1541.540 1.120 ;
  LAYER metal4 ;
  RECT 1538.000 0.000 1541.540 1.120 ;
  LAYER metal3 ;
  RECT 1538.000 0.000 1541.540 1.120 ;
  LAYER metal2 ;
  RECT 1538.000 0.000 1541.540 1.120 ;
  LAYER metal1 ;
  RECT 1538.000 0.000 1541.540 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1524.360 0.000 1527.900 1.120 ;
  LAYER metal4 ;
  RECT 1524.360 0.000 1527.900 1.120 ;
  LAYER metal3 ;
  RECT 1524.360 0.000 1527.900 1.120 ;
  LAYER metal2 ;
  RECT 1524.360 0.000 1527.900 1.120 ;
  LAYER metal1 ;
  RECT 1524.360 0.000 1527.900 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1511.340 0.000 1514.880 1.120 ;
  LAYER metal4 ;
  RECT 1511.340 0.000 1514.880 1.120 ;
  LAYER metal3 ;
  RECT 1511.340 0.000 1514.880 1.120 ;
  LAYER metal2 ;
  RECT 1511.340 0.000 1514.880 1.120 ;
  LAYER metal1 ;
  RECT 1511.340 0.000 1514.880 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1497.700 0.000 1501.240 1.120 ;
  LAYER metal4 ;
  RECT 1497.700 0.000 1501.240 1.120 ;
  LAYER metal3 ;
  RECT 1497.700 0.000 1501.240 1.120 ;
  LAYER metal2 ;
  RECT 1497.700 0.000 1501.240 1.120 ;
  LAYER metal1 ;
  RECT 1497.700 0.000 1501.240 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1484.060 0.000 1487.600 1.120 ;
  LAYER metal4 ;
  RECT 1484.060 0.000 1487.600 1.120 ;
  LAYER metal3 ;
  RECT 1484.060 0.000 1487.600 1.120 ;
  LAYER metal2 ;
  RECT 1484.060 0.000 1487.600 1.120 ;
  LAYER metal1 ;
  RECT 1484.060 0.000 1487.600 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1417.100 0.000 1420.640 1.120 ;
  LAYER metal4 ;
  RECT 1417.100 0.000 1420.640 1.120 ;
  LAYER metal3 ;
  RECT 1417.100 0.000 1420.640 1.120 ;
  LAYER metal2 ;
  RECT 1417.100 0.000 1420.640 1.120 ;
  LAYER metal1 ;
  RECT 1417.100 0.000 1420.640 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1403.460 0.000 1407.000 1.120 ;
  LAYER metal4 ;
  RECT 1403.460 0.000 1407.000 1.120 ;
  LAYER metal3 ;
  RECT 1403.460 0.000 1407.000 1.120 ;
  LAYER metal2 ;
  RECT 1403.460 0.000 1407.000 1.120 ;
  LAYER metal1 ;
  RECT 1403.460 0.000 1407.000 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1390.440 0.000 1393.980 1.120 ;
  LAYER metal4 ;
  RECT 1390.440 0.000 1393.980 1.120 ;
  LAYER metal3 ;
  RECT 1390.440 0.000 1393.980 1.120 ;
  LAYER metal2 ;
  RECT 1390.440 0.000 1393.980 1.120 ;
  LAYER metal1 ;
  RECT 1390.440 0.000 1393.980 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1376.800 0.000 1380.340 1.120 ;
  LAYER metal4 ;
  RECT 1376.800 0.000 1380.340 1.120 ;
  LAYER metal3 ;
  RECT 1376.800 0.000 1380.340 1.120 ;
  LAYER metal2 ;
  RECT 1376.800 0.000 1380.340 1.120 ;
  LAYER metal1 ;
  RECT 1376.800 0.000 1380.340 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1363.160 0.000 1366.700 1.120 ;
  LAYER metal4 ;
  RECT 1363.160 0.000 1366.700 1.120 ;
  LAYER metal3 ;
  RECT 1363.160 0.000 1366.700 1.120 ;
  LAYER metal2 ;
  RECT 1363.160 0.000 1366.700 1.120 ;
  LAYER metal1 ;
  RECT 1363.160 0.000 1366.700 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1350.140 0.000 1353.680 1.120 ;
  LAYER metal4 ;
  RECT 1350.140 0.000 1353.680 1.120 ;
  LAYER metal3 ;
  RECT 1350.140 0.000 1353.680 1.120 ;
  LAYER metal2 ;
  RECT 1350.140 0.000 1353.680 1.120 ;
  LAYER metal1 ;
  RECT 1350.140 0.000 1353.680 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1282.560 0.000 1286.100 1.120 ;
  LAYER metal4 ;
  RECT 1282.560 0.000 1286.100 1.120 ;
  LAYER metal3 ;
  RECT 1282.560 0.000 1286.100 1.120 ;
  LAYER metal2 ;
  RECT 1282.560 0.000 1286.100 1.120 ;
  LAYER metal1 ;
  RECT 1282.560 0.000 1286.100 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1268.920 0.000 1272.460 1.120 ;
  LAYER metal4 ;
  RECT 1268.920 0.000 1272.460 1.120 ;
  LAYER metal3 ;
  RECT 1268.920 0.000 1272.460 1.120 ;
  LAYER metal2 ;
  RECT 1268.920 0.000 1272.460 1.120 ;
  LAYER metal1 ;
  RECT 1268.920 0.000 1272.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1255.900 0.000 1259.440 1.120 ;
  LAYER metal4 ;
  RECT 1255.900 0.000 1259.440 1.120 ;
  LAYER metal3 ;
  RECT 1255.900 0.000 1259.440 1.120 ;
  LAYER metal2 ;
  RECT 1255.900 0.000 1259.440 1.120 ;
  LAYER metal1 ;
  RECT 1255.900 0.000 1259.440 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1242.260 0.000 1245.800 1.120 ;
  LAYER metal4 ;
  RECT 1242.260 0.000 1245.800 1.120 ;
  LAYER metal3 ;
  RECT 1242.260 0.000 1245.800 1.120 ;
  LAYER metal2 ;
  RECT 1242.260 0.000 1245.800 1.120 ;
  LAYER metal1 ;
  RECT 1242.260 0.000 1245.800 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1228.620 0.000 1232.160 1.120 ;
  LAYER metal4 ;
  RECT 1228.620 0.000 1232.160 1.120 ;
  LAYER metal3 ;
  RECT 1228.620 0.000 1232.160 1.120 ;
  LAYER metal2 ;
  RECT 1228.620 0.000 1232.160 1.120 ;
  LAYER metal1 ;
  RECT 1228.620 0.000 1232.160 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1215.600 0.000 1219.140 1.120 ;
  LAYER metal4 ;
  RECT 1215.600 0.000 1219.140 1.120 ;
  LAYER metal3 ;
  RECT 1215.600 0.000 1219.140 1.120 ;
  LAYER metal2 ;
  RECT 1215.600 0.000 1219.140 1.120 ;
  LAYER metal1 ;
  RECT 1215.600 0.000 1219.140 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1148.020 0.000 1151.560 1.120 ;
  LAYER metal4 ;
  RECT 1148.020 0.000 1151.560 1.120 ;
  LAYER metal3 ;
  RECT 1148.020 0.000 1151.560 1.120 ;
  LAYER metal2 ;
  RECT 1148.020 0.000 1151.560 1.120 ;
  LAYER metal1 ;
  RECT 1148.020 0.000 1151.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1135.000 0.000 1138.540 1.120 ;
  LAYER metal4 ;
  RECT 1135.000 0.000 1138.540 1.120 ;
  LAYER metal3 ;
  RECT 1135.000 0.000 1138.540 1.120 ;
  LAYER metal2 ;
  RECT 1135.000 0.000 1138.540 1.120 ;
  LAYER metal1 ;
  RECT 1135.000 0.000 1138.540 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1121.360 0.000 1124.900 1.120 ;
  LAYER metal4 ;
  RECT 1121.360 0.000 1124.900 1.120 ;
  LAYER metal3 ;
  RECT 1121.360 0.000 1124.900 1.120 ;
  LAYER metal2 ;
  RECT 1121.360 0.000 1124.900 1.120 ;
  LAYER metal1 ;
  RECT 1121.360 0.000 1124.900 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1107.720 0.000 1111.260 1.120 ;
  LAYER metal4 ;
  RECT 1107.720 0.000 1111.260 1.120 ;
  LAYER metal3 ;
  RECT 1107.720 0.000 1111.260 1.120 ;
  LAYER metal2 ;
  RECT 1107.720 0.000 1111.260 1.120 ;
  LAYER metal1 ;
  RECT 1107.720 0.000 1111.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1094.700 0.000 1098.240 1.120 ;
  LAYER metal4 ;
  RECT 1094.700 0.000 1098.240 1.120 ;
  LAYER metal3 ;
  RECT 1094.700 0.000 1098.240 1.120 ;
  LAYER metal2 ;
  RECT 1094.700 0.000 1098.240 1.120 ;
  LAYER metal1 ;
  RECT 1094.700 0.000 1098.240 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1081.060 0.000 1084.600 1.120 ;
  LAYER metal4 ;
  RECT 1081.060 0.000 1084.600 1.120 ;
  LAYER metal3 ;
  RECT 1081.060 0.000 1084.600 1.120 ;
  LAYER metal2 ;
  RECT 1081.060 0.000 1084.600 1.120 ;
  LAYER metal1 ;
  RECT 1081.060 0.000 1084.600 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1014.100 0.000 1017.640 1.120 ;
  LAYER metal4 ;
  RECT 1014.100 0.000 1017.640 1.120 ;
  LAYER metal3 ;
  RECT 1014.100 0.000 1017.640 1.120 ;
  LAYER metal2 ;
  RECT 1014.100 0.000 1017.640 1.120 ;
  LAYER metal1 ;
  RECT 1014.100 0.000 1017.640 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 1000.460 0.000 1004.000 1.120 ;
  LAYER metal4 ;
  RECT 1000.460 0.000 1004.000 1.120 ;
  LAYER metal3 ;
  RECT 1000.460 0.000 1004.000 1.120 ;
  LAYER metal2 ;
  RECT 1000.460 0.000 1004.000 1.120 ;
  LAYER metal1 ;
  RECT 1000.460 0.000 1004.000 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 986.820 0.000 990.360 1.120 ;
  LAYER metal4 ;
  RECT 986.820 0.000 990.360 1.120 ;
  LAYER metal3 ;
  RECT 986.820 0.000 990.360 1.120 ;
  LAYER metal2 ;
  RECT 986.820 0.000 990.360 1.120 ;
  LAYER metal1 ;
  RECT 986.820 0.000 990.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 973.800 0.000 977.340 1.120 ;
  LAYER metal4 ;
  RECT 973.800 0.000 977.340 1.120 ;
  LAYER metal3 ;
  RECT 973.800 0.000 977.340 1.120 ;
  LAYER metal2 ;
  RECT 973.800 0.000 977.340 1.120 ;
  LAYER metal1 ;
  RECT 973.800 0.000 977.340 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 960.160 0.000 963.700 1.120 ;
  LAYER metal4 ;
  RECT 960.160 0.000 963.700 1.120 ;
  LAYER metal3 ;
  RECT 960.160 0.000 963.700 1.120 ;
  LAYER metal2 ;
  RECT 960.160 0.000 963.700 1.120 ;
  LAYER metal1 ;
  RECT 960.160 0.000 963.700 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 946.520 0.000 950.060 1.120 ;
  LAYER metal4 ;
  RECT 946.520 0.000 950.060 1.120 ;
  LAYER metal3 ;
  RECT 946.520 0.000 950.060 1.120 ;
  LAYER metal2 ;
  RECT 946.520 0.000 950.060 1.120 ;
  LAYER metal1 ;
  RECT 946.520 0.000 950.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 879.560 0.000 883.100 1.120 ;
  LAYER metal4 ;
  RECT 879.560 0.000 883.100 1.120 ;
  LAYER metal3 ;
  RECT 879.560 0.000 883.100 1.120 ;
  LAYER metal2 ;
  RECT 879.560 0.000 883.100 1.120 ;
  LAYER metal1 ;
  RECT 879.560 0.000 883.100 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 865.920 0.000 869.460 1.120 ;
  LAYER metal4 ;
  RECT 865.920 0.000 869.460 1.120 ;
  LAYER metal3 ;
  RECT 865.920 0.000 869.460 1.120 ;
  LAYER metal2 ;
  RECT 865.920 0.000 869.460 1.120 ;
  LAYER metal1 ;
  RECT 865.920 0.000 869.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 852.280 0.000 855.820 1.120 ;
  LAYER metal4 ;
  RECT 852.280 0.000 855.820 1.120 ;
  LAYER metal3 ;
  RECT 852.280 0.000 855.820 1.120 ;
  LAYER metal2 ;
  RECT 852.280 0.000 855.820 1.120 ;
  LAYER metal1 ;
  RECT 852.280 0.000 855.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 839.260 0.000 842.800 1.120 ;
  LAYER metal4 ;
  RECT 839.260 0.000 842.800 1.120 ;
  LAYER metal3 ;
  RECT 839.260 0.000 842.800 1.120 ;
  LAYER metal2 ;
  RECT 839.260 0.000 842.800 1.120 ;
  LAYER metal1 ;
  RECT 839.260 0.000 842.800 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 825.620 0.000 829.160 1.120 ;
  LAYER metal4 ;
  RECT 825.620 0.000 829.160 1.120 ;
  LAYER metal3 ;
  RECT 825.620 0.000 829.160 1.120 ;
  LAYER metal2 ;
  RECT 825.620 0.000 829.160 1.120 ;
  LAYER metal1 ;
  RECT 825.620 0.000 829.160 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 811.980 0.000 815.520 1.120 ;
  LAYER metal4 ;
  RECT 811.980 0.000 815.520 1.120 ;
  LAYER metal3 ;
  RECT 811.980 0.000 815.520 1.120 ;
  LAYER metal2 ;
  RECT 811.980 0.000 815.520 1.120 ;
  LAYER metal1 ;
  RECT 811.980 0.000 815.520 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 745.020 0.000 748.560 1.120 ;
  LAYER metal4 ;
  RECT 745.020 0.000 748.560 1.120 ;
  LAYER metal3 ;
  RECT 745.020 0.000 748.560 1.120 ;
  LAYER metal2 ;
  RECT 745.020 0.000 748.560 1.120 ;
  LAYER metal1 ;
  RECT 745.020 0.000 748.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 731.380 0.000 734.920 1.120 ;
  LAYER metal4 ;
  RECT 731.380 0.000 734.920 1.120 ;
  LAYER metal3 ;
  RECT 731.380 0.000 734.920 1.120 ;
  LAYER metal2 ;
  RECT 731.380 0.000 734.920 1.120 ;
  LAYER metal1 ;
  RECT 731.380 0.000 734.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 718.360 0.000 721.900 1.120 ;
  LAYER metal4 ;
  RECT 718.360 0.000 721.900 1.120 ;
  LAYER metal3 ;
  RECT 718.360 0.000 721.900 1.120 ;
  LAYER metal2 ;
  RECT 718.360 0.000 721.900 1.120 ;
  LAYER metal1 ;
  RECT 718.360 0.000 721.900 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 704.720 0.000 708.260 1.120 ;
  LAYER metal4 ;
  RECT 704.720 0.000 708.260 1.120 ;
  LAYER metal3 ;
  RECT 704.720 0.000 708.260 1.120 ;
  LAYER metal2 ;
  RECT 704.720 0.000 708.260 1.120 ;
  LAYER metal1 ;
  RECT 704.720 0.000 708.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 691.080 0.000 694.620 1.120 ;
  LAYER metal4 ;
  RECT 691.080 0.000 694.620 1.120 ;
  LAYER metal3 ;
  RECT 691.080 0.000 694.620 1.120 ;
  LAYER metal2 ;
  RECT 691.080 0.000 694.620 1.120 ;
  LAYER metal1 ;
  RECT 691.080 0.000 694.620 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 678.060 0.000 681.600 1.120 ;
  LAYER metal4 ;
  RECT 678.060 0.000 681.600 1.120 ;
  LAYER metal3 ;
  RECT 678.060 0.000 681.600 1.120 ;
  LAYER metal2 ;
  RECT 678.060 0.000 681.600 1.120 ;
  LAYER metal1 ;
  RECT 678.060 0.000 681.600 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 610.480 0.000 614.020 1.120 ;
  LAYER metal4 ;
  RECT 610.480 0.000 614.020 1.120 ;
  LAYER metal3 ;
  RECT 610.480 0.000 614.020 1.120 ;
  LAYER metal2 ;
  RECT 610.480 0.000 614.020 1.120 ;
  LAYER metal1 ;
  RECT 610.480 0.000 614.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 597.460 0.000 601.000 1.120 ;
  LAYER metal4 ;
  RECT 597.460 0.000 601.000 1.120 ;
  LAYER metal3 ;
  RECT 597.460 0.000 601.000 1.120 ;
  LAYER metal2 ;
  RECT 597.460 0.000 601.000 1.120 ;
  LAYER metal1 ;
  RECT 597.460 0.000 601.000 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 583.820 0.000 587.360 1.120 ;
  LAYER metal4 ;
  RECT 583.820 0.000 587.360 1.120 ;
  LAYER metal3 ;
  RECT 583.820 0.000 587.360 1.120 ;
  LAYER metal2 ;
  RECT 583.820 0.000 587.360 1.120 ;
  LAYER metal1 ;
  RECT 583.820 0.000 587.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 570.180 0.000 573.720 1.120 ;
  LAYER metal4 ;
  RECT 570.180 0.000 573.720 1.120 ;
  LAYER metal3 ;
  RECT 570.180 0.000 573.720 1.120 ;
  LAYER metal2 ;
  RECT 570.180 0.000 573.720 1.120 ;
  LAYER metal1 ;
  RECT 570.180 0.000 573.720 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 557.160 0.000 560.700 1.120 ;
  LAYER metal4 ;
  RECT 557.160 0.000 560.700 1.120 ;
  LAYER metal3 ;
  RECT 557.160 0.000 560.700 1.120 ;
  LAYER metal2 ;
  RECT 557.160 0.000 560.700 1.120 ;
  LAYER metal1 ;
  RECT 557.160 0.000 560.700 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 543.520 0.000 547.060 1.120 ;
  LAYER metal4 ;
  RECT 543.520 0.000 547.060 1.120 ;
  LAYER metal3 ;
  RECT 543.520 0.000 547.060 1.120 ;
  LAYER metal2 ;
  RECT 543.520 0.000 547.060 1.120 ;
  LAYER metal1 ;
  RECT 543.520 0.000 547.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 475.940 0.000 479.480 1.120 ;
  LAYER metal4 ;
  RECT 475.940 0.000 479.480 1.120 ;
  LAYER metal3 ;
  RECT 475.940 0.000 479.480 1.120 ;
  LAYER metal2 ;
  RECT 475.940 0.000 479.480 1.120 ;
  LAYER metal1 ;
  RECT 475.940 0.000 479.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 462.920 0.000 466.460 1.120 ;
  LAYER metal4 ;
  RECT 462.920 0.000 466.460 1.120 ;
  LAYER metal3 ;
  RECT 462.920 0.000 466.460 1.120 ;
  LAYER metal2 ;
  RECT 462.920 0.000 466.460 1.120 ;
  LAYER metal1 ;
  RECT 462.920 0.000 466.460 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 449.280 0.000 452.820 1.120 ;
  LAYER metal4 ;
  RECT 449.280 0.000 452.820 1.120 ;
  LAYER metal3 ;
  RECT 449.280 0.000 452.820 1.120 ;
  LAYER metal2 ;
  RECT 449.280 0.000 452.820 1.120 ;
  LAYER metal1 ;
  RECT 449.280 0.000 452.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 435.640 0.000 439.180 1.120 ;
  LAYER metal4 ;
  RECT 435.640 0.000 439.180 1.120 ;
  LAYER metal3 ;
  RECT 435.640 0.000 439.180 1.120 ;
  LAYER metal2 ;
  RECT 435.640 0.000 439.180 1.120 ;
  LAYER metal1 ;
  RECT 435.640 0.000 439.180 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 422.620 0.000 426.160 1.120 ;
  LAYER metal4 ;
  RECT 422.620 0.000 426.160 1.120 ;
  LAYER metal3 ;
  RECT 422.620 0.000 426.160 1.120 ;
  LAYER metal2 ;
  RECT 422.620 0.000 426.160 1.120 ;
  LAYER metal1 ;
  RECT 422.620 0.000 426.160 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 408.980 0.000 412.520 1.120 ;
  LAYER metal4 ;
  RECT 408.980 0.000 412.520 1.120 ;
  LAYER metal3 ;
  RECT 408.980 0.000 412.520 1.120 ;
  LAYER metal2 ;
  RECT 408.980 0.000 412.520 1.120 ;
  LAYER metal1 ;
  RECT 408.980 0.000 412.520 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 342.020 0.000 345.560 1.120 ;
  LAYER metal4 ;
  RECT 342.020 0.000 345.560 1.120 ;
  LAYER metal3 ;
  RECT 342.020 0.000 345.560 1.120 ;
  LAYER metal2 ;
  RECT 342.020 0.000 345.560 1.120 ;
  LAYER metal1 ;
  RECT 342.020 0.000 345.560 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 328.380 0.000 331.920 1.120 ;
  LAYER metal4 ;
  RECT 328.380 0.000 331.920 1.120 ;
  LAYER metal3 ;
  RECT 328.380 0.000 331.920 1.120 ;
  LAYER metal2 ;
  RECT 328.380 0.000 331.920 1.120 ;
  LAYER metal1 ;
  RECT 328.380 0.000 331.920 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 314.740 0.000 318.280 1.120 ;
  LAYER metal4 ;
  RECT 314.740 0.000 318.280 1.120 ;
  LAYER metal3 ;
  RECT 314.740 0.000 318.280 1.120 ;
  LAYER metal2 ;
  RECT 314.740 0.000 318.280 1.120 ;
  LAYER metal1 ;
  RECT 314.740 0.000 318.280 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 301.720 0.000 305.260 1.120 ;
  LAYER metal4 ;
  RECT 301.720 0.000 305.260 1.120 ;
  LAYER metal3 ;
  RECT 301.720 0.000 305.260 1.120 ;
  LAYER metal2 ;
  RECT 301.720 0.000 305.260 1.120 ;
  LAYER metal1 ;
  RECT 301.720 0.000 305.260 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 288.080 0.000 291.620 1.120 ;
  LAYER metal4 ;
  RECT 288.080 0.000 291.620 1.120 ;
  LAYER metal3 ;
  RECT 288.080 0.000 291.620 1.120 ;
  LAYER metal2 ;
  RECT 288.080 0.000 291.620 1.120 ;
  LAYER metal1 ;
  RECT 288.080 0.000 291.620 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 274.440 0.000 277.980 1.120 ;
  LAYER metal4 ;
  RECT 274.440 0.000 277.980 1.120 ;
  LAYER metal3 ;
  RECT 274.440 0.000 277.980 1.120 ;
  LAYER metal2 ;
  RECT 274.440 0.000 277.980 1.120 ;
  LAYER metal1 ;
  RECT 274.440 0.000 277.980 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 207.480 0.000 211.020 1.120 ;
  LAYER metal4 ;
  RECT 207.480 0.000 211.020 1.120 ;
  LAYER metal3 ;
  RECT 207.480 0.000 211.020 1.120 ;
  LAYER metal2 ;
  RECT 207.480 0.000 211.020 1.120 ;
  LAYER metal1 ;
  RECT 207.480 0.000 211.020 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 193.840 0.000 197.380 1.120 ;
  LAYER metal4 ;
  RECT 193.840 0.000 197.380 1.120 ;
  LAYER metal3 ;
  RECT 193.840 0.000 197.380 1.120 ;
  LAYER metal2 ;
  RECT 193.840 0.000 197.380 1.120 ;
  LAYER metal1 ;
  RECT 193.840 0.000 197.380 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 180.820 0.000 184.360 1.120 ;
  LAYER metal4 ;
  RECT 180.820 0.000 184.360 1.120 ;
  LAYER metal3 ;
  RECT 180.820 0.000 184.360 1.120 ;
  LAYER metal2 ;
  RECT 180.820 0.000 184.360 1.120 ;
  LAYER metal1 ;
  RECT 180.820 0.000 184.360 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 167.180 0.000 170.720 1.120 ;
  LAYER metal4 ;
  RECT 167.180 0.000 170.720 1.120 ;
  LAYER metal3 ;
  RECT 167.180 0.000 170.720 1.120 ;
  LAYER metal2 ;
  RECT 167.180 0.000 170.720 1.120 ;
  LAYER metal1 ;
  RECT 167.180 0.000 170.720 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 153.540 0.000 157.080 1.120 ;
  LAYER metal4 ;
  RECT 153.540 0.000 157.080 1.120 ;
  LAYER metal3 ;
  RECT 153.540 0.000 157.080 1.120 ;
  LAYER metal2 ;
  RECT 153.540 0.000 157.080 1.120 ;
  LAYER metal1 ;
  RECT 153.540 0.000 157.080 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 140.520 0.000 144.060 1.120 ;
  LAYER metal4 ;
  RECT 140.520 0.000 144.060 1.120 ;
  LAYER metal3 ;
  RECT 140.520 0.000 144.060 1.120 ;
  LAYER metal2 ;
  RECT 140.520 0.000 144.060 1.120 ;
  LAYER metal1 ;
  RECT 140.520 0.000 144.060 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 72.940 0.000 76.480 1.120 ;
  LAYER metal4 ;
  RECT 72.940 0.000 76.480 1.120 ;
  LAYER metal3 ;
  RECT 72.940 0.000 76.480 1.120 ;
  LAYER metal2 ;
  RECT 72.940 0.000 76.480 1.120 ;
  LAYER metal1 ;
  RECT 72.940 0.000 76.480 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 59.300 0.000 62.840 1.120 ;
  LAYER metal4 ;
  RECT 59.300 0.000 62.840 1.120 ;
  LAYER metal3 ;
  RECT 59.300 0.000 62.840 1.120 ;
  LAYER metal2 ;
  RECT 59.300 0.000 62.840 1.120 ;
  LAYER metal1 ;
  RECT 59.300 0.000 62.840 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 46.280 0.000 49.820 1.120 ;
  LAYER metal4 ;
  RECT 46.280 0.000 49.820 1.120 ;
  LAYER metal3 ;
  RECT 46.280 0.000 49.820 1.120 ;
  LAYER metal2 ;
  RECT 46.280 0.000 49.820 1.120 ;
  LAYER metal1 ;
  RECT 46.280 0.000 49.820 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 32.640 0.000 36.180 1.120 ;
  LAYER metal4 ;
  RECT 32.640 0.000 36.180 1.120 ;
  LAYER metal3 ;
  RECT 32.640 0.000 36.180 1.120 ;
  LAYER metal2 ;
  RECT 32.640 0.000 36.180 1.120 ;
  LAYER metal1 ;
  RECT 32.640 0.000 36.180 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 19.000 0.000 22.540 1.120 ;
  LAYER metal4 ;
  RECT 19.000 0.000 22.540 1.120 ;
  LAYER metal3 ;
  RECT 19.000 0.000 22.540 1.120 ;
  LAYER metal2 ;
  RECT 19.000 0.000 22.540 1.120 ;
  LAYER metal1 ;
  RECT 19.000 0.000 22.540 1.120 ;
 END
 PORT
  LAYER metal5 ;
  RECT 7.220 0.000 10.760 1.120 ;
  LAYER metal4 ;
  RECT 7.220 0.000 10.760 1.120 ;
  LAYER metal3 ;
  RECT 7.220 0.000 10.760 1.120 ;
  LAYER metal2 ;
  RECT 7.220 0.000 10.760 1.120 ;
  LAYER metal1 ;
  RECT 7.220 0.000 10.760 1.120 ;
 END
END VCC
PIN DIB127
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3548.940 208.880 3550.060 210.000 ;
  LAYER metal4 ;
  RECT 3548.940 208.880 3550.060 210.000 ;
  LAYER metal3 ;
  RECT 3548.940 208.880 3550.060 210.000 ;
  LAYER metal2 ;
  RECT 3548.940 208.880 3550.060 210.000 ;
  LAYER metal1 ;
  RECT 3548.940 208.880 3550.060 210.000 ;
 END
END DIB127
PIN DOB127
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3535.300 208.880 3536.420 210.000 ;
  LAYER metal4 ;
  RECT 3535.300 208.880 3536.420 210.000 ;
  LAYER metal3 ;
  RECT 3535.300 208.880 3536.420 210.000 ;
  LAYER metal2 ;
  RECT 3535.300 208.880 3536.420 210.000 ;
  LAYER metal1 ;
  RECT 3535.300 208.880 3536.420 210.000 ;
 END
END DOB127
PIN DIB126
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3522.280 208.880 3523.400 210.000 ;
  LAYER metal4 ;
  RECT 3522.280 208.880 3523.400 210.000 ;
  LAYER metal3 ;
  RECT 3522.280 208.880 3523.400 210.000 ;
  LAYER metal2 ;
  RECT 3522.280 208.880 3523.400 210.000 ;
  LAYER metal1 ;
  RECT 3522.280 208.880 3523.400 210.000 ;
 END
END DIB126
PIN DOB126
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3508.640 208.880 3509.760 210.000 ;
  LAYER metal4 ;
  RECT 3508.640 208.880 3509.760 210.000 ;
  LAYER metal3 ;
  RECT 3508.640 208.880 3509.760 210.000 ;
  LAYER metal2 ;
  RECT 3508.640 208.880 3509.760 210.000 ;
  LAYER metal1 ;
  RECT 3508.640 208.880 3509.760 210.000 ;
 END
END DOB126
PIN DIB125
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3495.000 208.880 3496.120 210.000 ;
  LAYER metal4 ;
  RECT 3495.000 208.880 3496.120 210.000 ;
  LAYER metal3 ;
  RECT 3495.000 208.880 3496.120 210.000 ;
  LAYER metal2 ;
  RECT 3495.000 208.880 3496.120 210.000 ;
  LAYER metal1 ;
  RECT 3495.000 208.880 3496.120 210.000 ;
 END
END DIB125
PIN DOB125
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3481.980 208.880 3483.100 210.000 ;
  LAYER metal4 ;
  RECT 3481.980 208.880 3483.100 210.000 ;
  LAYER metal3 ;
  RECT 3481.980 208.880 3483.100 210.000 ;
  LAYER metal2 ;
  RECT 3481.980 208.880 3483.100 210.000 ;
  LAYER metal1 ;
  RECT 3481.980 208.880 3483.100 210.000 ;
 END
END DOB125
PIN DIB124
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3468.340 208.880 3469.460 210.000 ;
  LAYER metal4 ;
  RECT 3468.340 208.880 3469.460 210.000 ;
  LAYER metal3 ;
  RECT 3468.340 208.880 3469.460 210.000 ;
  LAYER metal2 ;
  RECT 3468.340 208.880 3469.460 210.000 ;
  LAYER metal1 ;
  RECT 3468.340 208.880 3469.460 210.000 ;
 END
END DIB124
PIN DOB124
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3454.700 208.880 3455.820 210.000 ;
  LAYER metal4 ;
  RECT 3454.700 208.880 3455.820 210.000 ;
  LAYER metal3 ;
  RECT 3454.700 208.880 3455.820 210.000 ;
  LAYER metal2 ;
  RECT 3454.700 208.880 3455.820 210.000 ;
  LAYER metal1 ;
  RECT 3454.700 208.880 3455.820 210.000 ;
 END
END DOB124
PIN DIB123
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3441.060 208.880 3442.180 210.000 ;
  LAYER metal4 ;
  RECT 3441.060 208.880 3442.180 210.000 ;
  LAYER metal3 ;
  RECT 3441.060 208.880 3442.180 210.000 ;
  LAYER metal2 ;
  RECT 3441.060 208.880 3442.180 210.000 ;
  LAYER metal1 ;
  RECT 3441.060 208.880 3442.180 210.000 ;
 END
END DIB123
PIN DOB123
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3428.040 208.880 3429.160 210.000 ;
  LAYER metal4 ;
  RECT 3428.040 208.880 3429.160 210.000 ;
  LAYER metal3 ;
  RECT 3428.040 208.880 3429.160 210.000 ;
  LAYER metal2 ;
  RECT 3428.040 208.880 3429.160 210.000 ;
  LAYER metal1 ;
  RECT 3428.040 208.880 3429.160 210.000 ;
 END
END DOB123
PIN DIB122
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3414.400 208.880 3415.520 210.000 ;
  LAYER metal4 ;
  RECT 3414.400 208.880 3415.520 210.000 ;
  LAYER metal3 ;
  RECT 3414.400 208.880 3415.520 210.000 ;
  LAYER metal2 ;
  RECT 3414.400 208.880 3415.520 210.000 ;
  LAYER metal1 ;
  RECT 3414.400 208.880 3415.520 210.000 ;
 END
END DIB122
PIN DOB122
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3400.760 208.880 3401.880 210.000 ;
  LAYER metal4 ;
  RECT 3400.760 208.880 3401.880 210.000 ;
  LAYER metal3 ;
  RECT 3400.760 208.880 3401.880 210.000 ;
  LAYER metal2 ;
  RECT 3400.760 208.880 3401.880 210.000 ;
  LAYER metal1 ;
  RECT 3400.760 208.880 3401.880 210.000 ;
 END
END DOB122
PIN DIB121
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3387.740 208.880 3388.860 210.000 ;
  LAYER metal4 ;
  RECT 3387.740 208.880 3388.860 210.000 ;
  LAYER metal3 ;
  RECT 3387.740 208.880 3388.860 210.000 ;
  LAYER metal2 ;
  RECT 3387.740 208.880 3388.860 210.000 ;
  LAYER metal1 ;
  RECT 3387.740 208.880 3388.860 210.000 ;
 END
END DIB121
PIN DOB121
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3374.100 208.880 3375.220 210.000 ;
  LAYER metal4 ;
  RECT 3374.100 208.880 3375.220 210.000 ;
  LAYER metal3 ;
  RECT 3374.100 208.880 3375.220 210.000 ;
  LAYER metal2 ;
  RECT 3374.100 208.880 3375.220 210.000 ;
  LAYER metal1 ;
  RECT 3374.100 208.880 3375.220 210.000 ;
 END
END DOB121
PIN DIB120
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3360.460 208.880 3361.580 210.000 ;
  LAYER metal4 ;
  RECT 3360.460 208.880 3361.580 210.000 ;
  LAYER metal3 ;
  RECT 3360.460 208.880 3361.580 210.000 ;
  LAYER metal2 ;
  RECT 3360.460 208.880 3361.580 210.000 ;
  LAYER metal1 ;
  RECT 3360.460 208.880 3361.580 210.000 ;
 END
END DIB120
PIN DOB120
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3347.440 208.880 3348.560 210.000 ;
  LAYER metal4 ;
  RECT 3347.440 208.880 3348.560 210.000 ;
  LAYER metal3 ;
  RECT 3347.440 208.880 3348.560 210.000 ;
  LAYER metal2 ;
  RECT 3347.440 208.880 3348.560 210.000 ;
  LAYER metal1 ;
  RECT 3347.440 208.880 3348.560 210.000 ;
 END
END DOB120
PIN DIB119
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3333.800 208.880 3334.920 210.000 ;
  LAYER metal4 ;
  RECT 3333.800 208.880 3334.920 210.000 ;
  LAYER metal3 ;
  RECT 3333.800 208.880 3334.920 210.000 ;
  LAYER metal2 ;
  RECT 3333.800 208.880 3334.920 210.000 ;
  LAYER metal1 ;
  RECT 3333.800 208.880 3334.920 210.000 ;
 END
END DIB119
PIN DOB119
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3320.160 208.880 3321.280 210.000 ;
  LAYER metal4 ;
  RECT 3320.160 208.880 3321.280 210.000 ;
  LAYER metal3 ;
  RECT 3320.160 208.880 3321.280 210.000 ;
  LAYER metal2 ;
  RECT 3320.160 208.880 3321.280 210.000 ;
  LAYER metal1 ;
  RECT 3320.160 208.880 3321.280 210.000 ;
 END
END DOB119
PIN DIB118
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3307.140 208.880 3308.260 210.000 ;
  LAYER metal4 ;
  RECT 3307.140 208.880 3308.260 210.000 ;
  LAYER metal3 ;
  RECT 3307.140 208.880 3308.260 210.000 ;
  LAYER metal2 ;
  RECT 3307.140 208.880 3308.260 210.000 ;
  LAYER metal1 ;
  RECT 3307.140 208.880 3308.260 210.000 ;
 END
END DIB118
PIN DOB118
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3293.500 208.880 3294.620 210.000 ;
  LAYER metal4 ;
  RECT 3293.500 208.880 3294.620 210.000 ;
  LAYER metal3 ;
  RECT 3293.500 208.880 3294.620 210.000 ;
  LAYER metal2 ;
  RECT 3293.500 208.880 3294.620 210.000 ;
  LAYER metal1 ;
  RECT 3293.500 208.880 3294.620 210.000 ;
 END
END DOB118
PIN DIB117
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3279.860 208.880 3280.980 210.000 ;
  LAYER metal4 ;
  RECT 3279.860 208.880 3280.980 210.000 ;
  LAYER metal3 ;
  RECT 3279.860 208.880 3280.980 210.000 ;
  LAYER metal2 ;
  RECT 3279.860 208.880 3280.980 210.000 ;
  LAYER metal1 ;
  RECT 3279.860 208.880 3280.980 210.000 ;
 END
END DIB117
PIN DOB117
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3266.840 208.880 3267.960 210.000 ;
  LAYER metal4 ;
  RECT 3266.840 208.880 3267.960 210.000 ;
  LAYER metal3 ;
  RECT 3266.840 208.880 3267.960 210.000 ;
  LAYER metal2 ;
  RECT 3266.840 208.880 3267.960 210.000 ;
  LAYER metal1 ;
  RECT 3266.840 208.880 3267.960 210.000 ;
 END
END DOB117
PIN DIB116
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3253.200 208.880 3254.320 210.000 ;
  LAYER metal4 ;
  RECT 3253.200 208.880 3254.320 210.000 ;
  LAYER metal3 ;
  RECT 3253.200 208.880 3254.320 210.000 ;
  LAYER metal2 ;
  RECT 3253.200 208.880 3254.320 210.000 ;
  LAYER metal1 ;
  RECT 3253.200 208.880 3254.320 210.000 ;
 END
END DIB116
PIN DOB116
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3239.560 208.880 3240.680 210.000 ;
  LAYER metal4 ;
  RECT 3239.560 208.880 3240.680 210.000 ;
  LAYER metal3 ;
  RECT 3239.560 208.880 3240.680 210.000 ;
  LAYER metal2 ;
  RECT 3239.560 208.880 3240.680 210.000 ;
  LAYER metal1 ;
  RECT 3239.560 208.880 3240.680 210.000 ;
 END
END DOB116
PIN DIB115
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3226.540 208.880 3227.660 210.000 ;
  LAYER metal4 ;
  RECT 3226.540 208.880 3227.660 210.000 ;
  LAYER metal3 ;
  RECT 3226.540 208.880 3227.660 210.000 ;
  LAYER metal2 ;
  RECT 3226.540 208.880 3227.660 210.000 ;
  LAYER metal1 ;
  RECT 3226.540 208.880 3227.660 210.000 ;
 END
END DIB115
PIN DOB115
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3212.900 208.880 3214.020 210.000 ;
  LAYER metal4 ;
  RECT 3212.900 208.880 3214.020 210.000 ;
  LAYER metal3 ;
  RECT 3212.900 208.880 3214.020 210.000 ;
  LAYER metal2 ;
  RECT 3212.900 208.880 3214.020 210.000 ;
  LAYER metal1 ;
  RECT 3212.900 208.880 3214.020 210.000 ;
 END
END DOB115
PIN DIB114
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3199.260 208.880 3200.380 210.000 ;
  LAYER metal4 ;
  RECT 3199.260 208.880 3200.380 210.000 ;
  LAYER metal3 ;
  RECT 3199.260 208.880 3200.380 210.000 ;
  LAYER metal2 ;
  RECT 3199.260 208.880 3200.380 210.000 ;
  LAYER metal1 ;
  RECT 3199.260 208.880 3200.380 210.000 ;
 END
END DIB114
PIN DOB114
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3186.240 208.880 3187.360 210.000 ;
  LAYER metal4 ;
  RECT 3186.240 208.880 3187.360 210.000 ;
  LAYER metal3 ;
  RECT 3186.240 208.880 3187.360 210.000 ;
  LAYER metal2 ;
  RECT 3186.240 208.880 3187.360 210.000 ;
  LAYER metal1 ;
  RECT 3186.240 208.880 3187.360 210.000 ;
 END
END DOB114
PIN DIB113
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3172.600 208.880 3173.720 210.000 ;
  LAYER metal4 ;
  RECT 3172.600 208.880 3173.720 210.000 ;
  LAYER metal3 ;
  RECT 3172.600 208.880 3173.720 210.000 ;
  LAYER metal2 ;
  RECT 3172.600 208.880 3173.720 210.000 ;
  LAYER metal1 ;
  RECT 3172.600 208.880 3173.720 210.000 ;
 END
END DIB113
PIN DOB113
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3158.960 208.880 3160.080 210.000 ;
  LAYER metal4 ;
  RECT 3158.960 208.880 3160.080 210.000 ;
  LAYER metal3 ;
  RECT 3158.960 208.880 3160.080 210.000 ;
  LAYER metal2 ;
  RECT 3158.960 208.880 3160.080 210.000 ;
  LAYER metal1 ;
  RECT 3158.960 208.880 3160.080 210.000 ;
 END
END DOB113
PIN DIB112
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3145.940 208.880 3147.060 210.000 ;
  LAYER metal4 ;
  RECT 3145.940 208.880 3147.060 210.000 ;
  LAYER metal3 ;
  RECT 3145.940 208.880 3147.060 210.000 ;
  LAYER metal2 ;
  RECT 3145.940 208.880 3147.060 210.000 ;
  LAYER metal1 ;
  RECT 3145.940 208.880 3147.060 210.000 ;
 END
END DIB112
PIN DOB112
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3132.300 208.880 3133.420 210.000 ;
  LAYER metal4 ;
  RECT 3132.300 208.880 3133.420 210.000 ;
  LAYER metal3 ;
  RECT 3132.300 208.880 3133.420 210.000 ;
  LAYER metal2 ;
  RECT 3132.300 208.880 3133.420 210.000 ;
  LAYER metal1 ;
  RECT 3132.300 208.880 3133.420 210.000 ;
 END
END DOB112
PIN DIB111
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3118.660 208.880 3119.780 210.000 ;
  LAYER metal4 ;
  RECT 3118.660 208.880 3119.780 210.000 ;
  LAYER metal3 ;
  RECT 3118.660 208.880 3119.780 210.000 ;
  LAYER metal2 ;
  RECT 3118.660 208.880 3119.780 210.000 ;
  LAYER metal1 ;
  RECT 3118.660 208.880 3119.780 210.000 ;
 END
END DIB111
PIN DOB111
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3105.640 208.880 3106.760 210.000 ;
  LAYER metal4 ;
  RECT 3105.640 208.880 3106.760 210.000 ;
  LAYER metal3 ;
  RECT 3105.640 208.880 3106.760 210.000 ;
  LAYER metal2 ;
  RECT 3105.640 208.880 3106.760 210.000 ;
  LAYER metal1 ;
  RECT 3105.640 208.880 3106.760 210.000 ;
 END
END DOB111
PIN DIB110
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3092.000 208.880 3093.120 210.000 ;
  LAYER metal4 ;
  RECT 3092.000 208.880 3093.120 210.000 ;
  LAYER metal3 ;
  RECT 3092.000 208.880 3093.120 210.000 ;
  LAYER metal2 ;
  RECT 3092.000 208.880 3093.120 210.000 ;
  LAYER metal1 ;
  RECT 3092.000 208.880 3093.120 210.000 ;
 END
END DIB110
PIN DOB110
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3078.360 208.880 3079.480 210.000 ;
  LAYER metal4 ;
  RECT 3078.360 208.880 3079.480 210.000 ;
  LAYER metal3 ;
  RECT 3078.360 208.880 3079.480 210.000 ;
  LAYER metal2 ;
  RECT 3078.360 208.880 3079.480 210.000 ;
  LAYER metal1 ;
  RECT 3078.360 208.880 3079.480 210.000 ;
 END
END DOB110
PIN DIB109
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3065.340 208.880 3066.460 210.000 ;
  LAYER metal4 ;
  RECT 3065.340 208.880 3066.460 210.000 ;
  LAYER metal3 ;
  RECT 3065.340 208.880 3066.460 210.000 ;
  LAYER metal2 ;
  RECT 3065.340 208.880 3066.460 210.000 ;
  LAYER metal1 ;
  RECT 3065.340 208.880 3066.460 210.000 ;
 END
END DIB109
PIN DOB109
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3051.700 208.880 3052.820 210.000 ;
  LAYER metal4 ;
  RECT 3051.700 208.880 3052.820 210.000 ;
  LAYER metal3 ;
  RECT 3051.700 208.880 3052.820 210.000 ;
  LAYER metal2 ;
  RECT 3051.700 208.880 3052.820 210.000 ;
  LAYER metal1 ;
  RECT 3051.700 208.880 3052.820 210.000 ;
 END
END DOB109
PIN DIB108
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3038.060 208.880 3039.180 210.000 ;
  LAYER metal4 ;
  RECT 3038.060 208.880 3039.180 210.000 ;
  LAYER metal3 ;
  RECT 3038.060 208.880 3039.180 210.000 ;
  LAYER metal2 ;
  RECT 3038.060 208.880 3039.180 210.000 ;
  LAYER metal1 ;
  RECT 3038.060 208.880 3039.180 210.000 ;
 END
END DIB108
PIN DOB108
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3024.420 208.880 3025.540 210.000 ;
  LAYER metal4 ;
  RECT 3024.420 208.880 3025.540 210.000 ;
  LAYER metal3 ;
  RECT 3024.420 208.880 3025.540 210.000 ;
  LAYER metal2 ;
  RECT 3024.420 208.880 3025.540 210.000 ;
  LAYER metal1 ;
  RECT 3024.420 208.880 3025.540 210.000 ;
 END
END DOB108
PIN DIB107
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3011.400 208.880 3012.520 210.000 ;
  LAYER metal4 ;
  RECT 3011.400 208.880 3012.520 210.000 ;
  LAYER metal3 ;
  RECT 3011.400 208.880 3012.520 210.000 ;
  LAYER metal2 ;
  RECT 3011.400 208.880 3012.520 210.000 ;
  LAYER metal1 ;
  RECT 3011.400 208.880 3012.520 210.000 ;
 END
END DIB107
PIN DOB107
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2997.760 208.880 2998.880 210.000 ;
  LAYER metal4 ;
  RECT 2997.760 208.880 2998.880 210.000 ;
  LAYER metal3 ;
  RECT 2997.760 208.880 2998.880 210.000 ;
  LAYER metal2 ;
  RECT 2997.760 208.880 2998.880 210.000 ;
  LAYER metal1 ;
  RECT 2997.760 208.880 2998.880 210.000 ;
 END
END DOB107
PIN DIB106
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2984.120 208.880 2985.240 210.000 ;
  LAYER metal4 ;
  RECT 2984.120 208.880 2985.240 210.000 ;
  LAYER metal3 ;
  RECT 2984.120 208.880 2985.240 210.000 ;
  LAYER metal2 ;
  RECT 2984.120 208.880 2985.240 210.000 ;
  LAYER metal1 ;
  RECT 2984.120 208.880 2985.240 210.000 ;
 END
END DIB106
PIN DOB106
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2971.100 208.880 2972.220 210.000 ;
  LAYER metal4 ;
  RECT 2971.100 208.880 2972.220 210.000 ;
  LAYER metal3 ;
  RECT 2971.100 208.880 2972.220 210.000 ;
  LAYER metal2 ;
  RECT 2971.100 208.880 2972.220 210.000 ;
  LAYER metal1 ;
  RECT 2971.100 208.880 2972.220 210.000 ;
 END
END DOB106
PIN DIB105
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2957.460 208.880 2958.580 210.000 ;
  LAYER metal4 ;
  RECT 2957.460 208.880 2958.580 210.000 ;
  LAYER metal3 ;
  RECT 2957.460 208.880 2958.580 210.000 ;
  LAYER metal2 ;
  RECT 2957.460 208.880 2958.580 210.000 ;
  LAYER metal1 ;
  RECT 2957.460 208.880 2958.580 210.000 ;
 END
END DIB105
PIN DOB105
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2943.820 208.880 2944.940 210.000 ;
  LAYER metal4 ;
  RECT 2943.820 208.880 2944.940 210.000 ;
  LAYER metal3 ;
  RECT 2943.820 208.880 2944.940 210.000 ;
  LAYER metal2 ;
  RECT 2943.820 208.880 2944.940 210.000 ;
  LAYER metal1 ;
  RECT 2943.820 208.880 2944.940 210.000 ;
 END
END DOB105
PIN DIB104
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2930.800 208.880 2931.920 210.000 ;
  LAYER metal4 ;
  RECT 2930.800 208.880 2931.920 210.000 ;
  LAYER metal3 ;
  RECT 2930.800 208.880 2931.920 210.000 ;
  LAYER metal2 ;
  RECT 2930.800 208.880 2931.920 210.000 ;
  LAYER metal1 ;
  RECT 2930.800 208.880 2931.920 210.000 ;
 END
END DIB104
PIN DOB104
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2917.160 208.880 2918.280 210.000 ;
  LAYER metal4 ;
  RECT 2917.160 208.880 2918.280 210.000 ;
  LAYER metal3 ;
  RECT 2917.160 208.880 2918.280 210.000 ;
  LAYER metal2 ;
  RECT 2917.160 208.880 2918.280 210.000 ;
  LAYER metal1 ;
  RECT 2917.160 208.880 2918.280 210.000 ;
 END
END DOB104
PIN DIB103
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2903.520 208.880 2904.640 210.000 ;
  LAYER metal4 ;
  RECT 2903.520 208.880 2904.640 210.000 ;
  LAYER metal3 ;
  RECT 2903.520 208.880 2904.640 210.000 ;
  LAYER metal2 ;
  RECT 2903.520 208.880 2904.640 210.000 ;
  LAYER metal1 ;
  RECT 2903.520 208.880 2904.640 210.000 ;
 END
END DIB103
PIN DOB103
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2890.500 208.880 2891.620 210.000 ;
  LAYER metal4 ;
  RECT 2890.500 208.880 2891.620 210.000 ;
  LAYER metal3 ;
  RECT 2890.500 208.880 2891.620 210.000 ;
  LAYER metal2 ;
  RECT 2890.500 208.880 2891.620 210.000 ;
  LAYER metal1 ;
  RECT 2890.500 208.880 2891.620 210.000 ;
 END
END DOB103
PIN DIB102
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2876.860 208.880 2877.980 210.000 ;
  LAYER metal4 ;
  RECT 2876.860 208.880 2877.980 210.000 ;
  LAYER metal3 ;
  RECT 2876.860 208.880 2877.980 210.000 ;
  LAYER metal2 ;
  RECT 2876.860 208.880 2877.980 210.000 ;
  LAYER metal1 ;
  RECT 2876.860 208.880 2877.980 210.000 ;
 END
END DIB102
PIN DOB102
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2863.220 208.880 2864.340 210.000 ;
  LAYER metal4 ;
  RECT 2863.220 208.880 2864.340 210.000 ;
  LAYER metal3 ;
  RECT 2863.220 208.880 2864.340 210.000 ;
  LAYER metal2 ;
  RECT 2863.220 208.880 2864.340 210.000 ;
  LAYER metal1 ;
  RECT 2863.220 208.880 2864.340 210.000 ;
 END
END DOB102
PIN DIB101
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2850.200 208.880 2851.320 210.000 ;
  LAYER metal4 ;
  RECT 2850.200 208.880 2851.320 210.000 ;
  LAYER metal3 ;
  RECT 2850.200 208.880 2851.320 210.000 ;
  LAYER metal2 ;
  RECT 2850.200 208.880 2851.320 210.000 ;
  LAYER metal1 ;
  RECT 2850.200 208.880 2851.320 210.000 ;
 END
END DIB101
PIN DOB101
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2836.560 208.880 2837.680 210.000 ;
  LAYER metal4 ;
  RECT 2836.560 208.880 2837.680 210.000 ;
  LAYER metal3 ;
  RECT 2836.560 208.880 2837.680 210.000 ;
  LAYER metal2 ;
  RECT 2836.560 208.880 2837.680 210.000 ;
  LAYER metal1 ;
  RECT 2836.560 208.880 2837.680 210.000 ;
 END
END DOB101
PIN DIB100
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2822.920 208.880 2824.040 210.000 ;
  LAYER metal4 ;
  RECT 2822.920 208.880 2824.040 210.000 ;
  LAYER metal3 ;
  RECT 2822.920 208.880 2824.040 210.000 ;
  LAYER metal2 ;
  RECT 2822.920 208.880 2824.040 210.000 ;
  LAYER metal1 ;
  RECT 2822.920 208.880 2824.040 210.000 ;
 END
END DIB100
PIN DOB100
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2809.900 208.880 2811.020 210.000 ;
  LAYER metal4 ;
  RECT 2809.900 208.880 2811.020 210.000 ;
  LAYER metal3 ;
  RECT 2809.900 208.880 2811.020 210.000 ;
  LAYER metal2 ;
  RECT 2809.900 208.880 2811.020 210.000 ;
  LAYER metal1 ;
  RECT 2809.900 208.880 2811.020 210.000 ;
 END
END DOB100
PIN DIB99
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2796.260 208.880 2797.380 210.000 ;
  LAYER metal4 ;
  RECT 2796.260 208.880 2797.380 210.000 ;
  LAYER metal3 ;
  RECT 2796.260 208.880 2797.380 210.000 ;
  LAYER metal2 ;
  RECT 2796.260 208.880 2797.380 210.000 ;
  LAYER metal1 ;
  RECT 2796.260 208.880 2797.380 210.000 ;
 END
END DIB99
PIN DOB99
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2782.620 208.880 2783.740 210.000 ;
  LAYER metal4 ;
  RECT 2782.620 208.880 2783.740 210.000 ;
  LAYER metal3 ;
  RECT 2782.620 208.880 2783.740 210.000 ;
  LAYER metal2 ;
  RECT 2782.620 208.880 2783.740 210.000 ;
  LAYER metal1 ;
  RECT 2782.620 208.880 2783.740 210.000 ;
 END
END DOB99
PIN DIB98
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2769.600 208.880 2770.720 210.000 ;
  LAYER metal4 ;
  RECT 2769.600 208.880 2770.720 210.000 ;
  LAYER metal3 ;
  RECT 2769.600 208.880 2770.720 210.000 ;
  LAYER metal2 ;
  RECT 2769.600 208.880 2770.720 210.000 ;
  LAYER metal1 ;
  RECT 2769.600 208.880 2770.720 210.000 ;
 END
END DIB98
PIN DOB98
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2755.960 208.880 2757.080 210.000 ;
  LAYER metal4 ;
  RECT 2755.960 208.880 2757.080 210.000 ;
  LAYER metal3 ;
  RECT 2755.960 208.880 2757.080 210.000 ;
  LAYER metal2 ;
  RECT 2755.960 208.880 2757.080 210.000 ;
  LAYER metal1 ;
  RECT 2755.960 208.880 2757.080 210.000 ;
 END
END DOB98
PIN DIB97
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2742.320 208.880 2743.440 210.000 ;
  LAYER metal4 ;
  RECT 2742.320 208.880 2743.440 210.000 ;
  LAYER metal3 ;
  RECT 2742.320 208.880 2743.440 210.000 ;
  LAYER metal2 ;
  RECT 2742.320 208.880 2743.440 210.000 ;
  LAYER metal1 ;
  RECT 2742.320 208.880 2743.440 210.000 ;
 END
END DIB97
PIN DOB97
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2729.300 208.880 2730.420 210.000 ;
  LAYER metal4 ;
  RECT 2729.300 208.880 2730.420 210.000 ;
  LAYER metal3 ;
  RECT 2729.300 208.880 2730.420 210.000 ;
  LAYER metal2 ;
  RECT 2729.300 208.880 2730.420 210.000 ;
  LAYER metal1 ;
  RECT 2729.300 208.880 2730.420 210.000 ;
 END
END DOB97
PIN DIB96
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2715.660 208.880 2716.780 210.000 ;
  LAYER metal4 ;
  RECT 2715.660 208.880 2716.780 210.000 ;
  LAYER metal3 ;
  RECT 2715.660 208.880 2716.780 210.000 ;
  LAYER metal2 ;
  RECT 2715.660 208.880 2716.780 210.000 ;
  LAYER metal1 ;
  RECT 2715.660 208.880 2716.780 210.000 ;
 END
END DIB96
PIN DOB96
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2702.020 208.880 2703.140 210.000 ;
  LAYER metal4 ;
  RECT 2702.020 208.880 2703.140 210.000 ;
  LAYER metal3 ;
  RECT 2702.020 208.880 2703.140 210.000 ;
  LAYER metal2 ;
  RECT 2702.020 208.880 2703.140 210.000 ;
  LAYER metal1 ;
  RECT 2702.020 208.880 2703.140 210.000 ;
 END
END DOB96
PIN DIB95
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2689.000 208.880 2690.120 210.000 ;
  LAYER metal4 ;
  RECT 2689.000 208.880 2690.120 210.000 ;
  LAYER metal3 ;
  RECT 2689.000 208.880 2690.120 210.000 ;
  LAYER metal2 ;
  RECT 2689.000 208.880 2690.120 210.000 ;
  LAYER metal1 ;
  RECT 2689.000 208.880 2690.120 210.000 ;
 END
END DIB95
PIN DOB95
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2675.360 208.880 2676.480 210.000 ;
  LAYER metal4 ;
  RECT 2675.360 208.880 2676.480 210.000 ;
  LAYER metal3 ;
  RECT 2675.360 208.880 2676.480 210.000 ;
  LAYER metal2 ;
  RECT 2675.360 208.880 2676.480 210.000 ;
  LAYER metal1 ;
  RECT 2675.360 208.880 2676.480 210.000 ;
 END
END DOB95
PIN DIB94
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2661.720 208.880 2662.840 210.000 ;
  LAYER metal4 ;
  RECT 2661.720 208.880 2662.840 210.000 ;
  LAYER metal3 ;
  RECT 2661.720 208.880 2662.840 210.000 ;
  LAYER metal2 ;
  RECT 2661.720 208.880 2662.840 210.000 ;
  LAYER metal1 ;
  RECT 2661.720 208.880 2662.840 210.000 ;
 END
END DIB94
PIN DOB94
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2648.700 208.880 2649.820 210.000 ;
  LAYER metal4 ;
  RECT 2648.700 208.880 2649.820 210.000 ;
  LAYER metal3 ;
  RECT 2648.700 208.880 2649.820 210.000 ;
  LAYER metal2 ;
  RECT 2648.700 208.880 2649.820 210.000 ;
  LAYER metal1 ;
  RECT 2648.700 208.880 2649.820 210.000 ;
 END
END DOB94
PIN DIB93
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2635.060 208.880 2636.180 210.000 ;
  LAYER metal4 ;
  RECT 2635.060 208.880 2636.180 210.000 ;
  LAYER metal3 ;
  RECT 2635.060 208.880 2636.180 210.000 ;
  LAYER metal2 ;
  RECT 2635.060 208.880 2636.180 210.000 ;
  LAYER metal1 ;
  RECT 2635.060 208.880 2636.180 210.000 ;
 END
END DIB93
PIN DOB93
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2621.420 208.880 2622.540 210.000 ;
  LAYER metal4 ;
  RECT 2621.420 208.880 2622.540 210.000 ;
  LAYER metal3 ;
  RECT 2621.420 208.880 2622.540 210.000 ;
  LAYER metal2 ;
  RECT 2621.420 208.880 2622.540 210.000 ;
  LAYER metal1 ;
  RECT 2621.420 208.880 2622.540 210.000 ;
 END
END DOB93
PIN DIB92
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2607.780 208.880 2608.900 210.000 ;
  LAYER metal4 ;
  RECT 2607.780 208.880 2608.900 210.000 ;
  LAYER metal3 ;
  RECT 2607.780 208.880 2608.900 210.000 ;
  LAYER metal2 ;
  RECT 2607.780 208.880 2608.900 210.000 ;
  LAYER metal1 ;
  RECT 2607.780 208.880 2608.900 210.000 ;
 END
END DIB92
PIN DOB92
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2594.760 208.880 2595.880 210.000 ;
  LAYER metal4 ;
  RECT 2594.760 208.880 2595.880 210.000 ;
  LAYER metal3 ;
  RECT 2594.760 208.880 2595.880 210.000 ;
  LAYER metal2 ;
  RECT 2594.760 208.880 2595.880 210.000 ;
  LAYER metal1 ;
  RECT 2594.760 208.880 2595.880 210.000 ;
 END
END DOB92
PIN DIB91
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2581.120 208.880 2582.240 210.000 ;
  LAYER metal4 ;
  RECT 2581.120 208.880 2582.240 210.000 ;
  LAYER metal3 ;
  RECT 2581.120 208.880 2582.240 210.000 ;
  LAYER metal2 ;
  RECT 2581.120 208.880 2582.240 210.000 ;
  LAYER metal1 ;
  RECT 2581.120 208.880 2582.240 210.000 ;
 END
END DIB91
PIN DOB91
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2567.480 208.880 2568.600 210.000 ;
  LAYER metal4 ;
  RECT 2567.480 208.880 2568.600 210.000 ;
  LAYER metal3 ;
  RECT 2567.480 208.880 2568.600 210.000 ;
  LAYER metal2 ;
  RECT 2567.480 208.880 2568.600 210.000 ;
  LAYER metal1 ;
  RECT 2567.480 208.880 2568.600 210.000 ;
 END
END DOB91
PIN DIB90
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2554.460 208.880 2555.580 210.000 ;
  LAYER metal4 ;
  RECT 2554.460 208.880 2555.580 210.000 ;
  LAYER metal3 ;
  RECT 2554.460 208.880 2555.580 210.000 ;
  LAYER metal2 ;
  RECT 2554.460 208.880 2555.580 210.000 ;
  LAYER metal1 ;
  RECT 2554.460 208.880 2555.580 210.000 ;
 END
END DIB90
PIN DOB90
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2540.820 208.880 2541.940 210.000 ;
  LAYER metal4 ;
  RECT 2540.820 208.880 2541.940 210.000 ;
  LAYER metal3 ;
  RECT 2540.820 208.880 2541.940 210.000 ;
  LAYER metal2 ;
  RECT 2540.820 208.880 2541.940 210.000 ;
  LAYER metal1 ;
  RECT 2540.820 208.880 2541.940 210.000 ;
 END
END DOB90
PIN DIB89
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2527.180 208.880 2528.300 210.000 ;
  LAYER metal4 ;
  RECT 2527.180 208.880 2528.300 210.000 ;
  LAYER metal3 ;
  RECT 2527.180 208.880 2528.300 210.000 ;
  LAYER metal2 ;
  RECT 2527.180 208.880 2528.300 210.000 ;
  LAYER metal1 ;
  RECT 2527.180 208.880 2528.300 210.000 ;
 END
END DIB89
PIN DOB89
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2514.160 208.880 2515.280 210.000 ;
  LAYER metal4 ;
  RECT 2514.160 208.880 2515.280 210.000 ;
  LAYER metal3 ;
  RECT 2514.160 208.880 2515.280 210.000 ;
  LAYER metal2 ;
  RECT 2514.160 208.880 2515.280 210.000 ;
  LAYER metal1 ;
  RECT 2514.160 208.880 2515.280 210.000 ;
 END
END DOB89
PIN DIB88
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2500.520 208.880 2501.640 210.000 ;
  LAYER metal4 ;
  RECT 2500.520 208.880 2501.640 210.000 ;
  LAYER metal3 ;
  RECT 2500.520 208.880 2501.640 210.000 ;
  LAYER metal2 ;
  RECT 2500.520 208.880 2501.640 210.000 ;
  LAYER metal1 ;
  RECT 2500.520 208.880 2501.640 210.000 ;
 END
END DIB88
PIN DOB88
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2486.880 208.880 2488.000 210.000 ;
  LAYER metal4 ;
  RECT 2486.880 208.880 2488.000 210.000 ;
  LAYER metal3 ;
  RECT 2486.880 208.880 2488.000 210.000 ;
  LAYER metal2 ;
  RECT 2486.880 208.880 2488.000 210.000 ;
  LAYER metal1 ;
  RECT 2486.880 208.880 2488.000 210.000 ;
 END
END DOB88
PIN DIB87
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2473.860 208.880 2474.980 210.000 ;
  LAYER metal4 ;
  RECT 2473.860 208.880 2474.980 210.000 ;
  LAYER metal3 ;
  RECT 2473.860 208.880 2474.980 210.000 ;
  LAYER metal2 ;
  RECT 2473.860 208.880 2474.980 210.000 ;
  LAYER metal1 ;
  RECT 2473.860 208.880 2474.980 210.000 ;
 END
END DIB87
PIN DOB87
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2460.220 208.880 2461.340 210.000 ;
  LAYER metal4 ;
  RECT 2460.220 208.880 2461.340 210.000 ;
  LAYER metal3 ;
  RECT 2460.220 208.880 2461.340 210.000 ;
  LAYER metal2 ;
  RECT 2460.220 208.880 2461.340 210.000 ;
  LAYER metal1 ;
  RECT 2460.220 208.880 2461.340 210.000 ;
 END
END DOB87
PIN DIB86
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2446.580 208.880 2447.700 210.000 ;
  LAYER metal4 ;
  RECT 2446.580 208.880 2447.700 210.000 ;
  LAYER metal3 ;
  RECT 2446.580 208.880 2447.700 210.000 ;
  LAYER metal2 ;
  RECT 2446.580 208.880 2447.700 210.000 ;
  LAYER metal1 ;
  RECT 2446.580 208.880 2447.700 210.000 ;
 END
END DIB86
PIN DOB86
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2433.560 208.880 2434.680 210.000 ;
  LAYER metal4 ;
  RECT 2433.560 208.880 2434.680 210.000 ;
  LAYER metal3 ;
  RECT 2433.560 208.880 2434.680 210.000 ;
  LAYER metal2 ;
  RECT 2433.560 208.880 2434.680 210.000 ;
  LAYER metal1 ;
  RECT 2433.560 208.880 2434.680 210.000 ;
 END
END DOB86
PIN DIB85
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2419.920 208.880 2421.040 210.000 ;
  LAYER metal4 ;
  RECT 2419.920 208.880 2421.040 210.000 ;
  LAYER metal3 ;
  RECT 2419.920 208.880 2421.040 210.000 ;
  LAYER metal2 ;
  RECT 2419.920 208.880 2421.040 210.000 ;
  LAYER metal1 ;
  RECT 2419.920 208.880 2421.040 210.000 ;
 END
END DIB85
PIN DOB85
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2406.280 208.880 2407.400 210.000 ;
  LAYER metal4 ;
  RECT 2406.280 208.880 2407.400 210.000 ;
  LAYER metal3 ;
  RECT 2406.280 208.880 2407.400 210.000 ;
  LAYER metal2 ;
  RECT 2406.280 208.880 2407.400 210.000 ;
  LAYER metal1 ;
  RECT 2406.280 208.880 2407.400 210.000 ;
 END
END DOB85
PIN DIB84
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2393.260 208.880 2394.380 210.000 ;
  LAYER metal4 ;
  RECT 2393.260 208.880 2394.380 210.000 ;
  LAYER metal3 ;
  RECT 2393.260 208.880 2394.380 210.000 ;
  LAYER metal2 ;
  RECT 2393.260 208.880 2394.380 210.000 ;
  LAYER metal1 ;
  RECT 2393.260 208.880 2394.380 210.000 ;
 END
END DIB84
PIN DOB84
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2379.620 208.880 2380.740 210.000 ;
  LAYER metal4 ;
  RECT 2379.620 208.880 2380.740 210.000 ;
  LAYER metal3 ;
  RECT 2379.620 208.880 2380.740 210.000 ;
  LAYER metal2 ;
  RECT 2379.620 208.880 2380.740 210.000 ;
  LAYER metal1 ;
  RECT 2379.620 208.880 2380.740 210.000 ;
 END
END DOB84
PIN DIB83
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2365.980 208.880 2367.100 210.000 ;
  LAYER metal4 ;
  RECT 2365.980 208.880 2367.100 210.000 ;
  LAYER metal3 ;
  RECT 2365.980 208.880 2367.100 210.000 ;
  LAYER metal2 ;
  RECT 2365.980 208.880 2367.100 210.000 ;
  LAYER metal1 ;
  RECT 2365.980 208.880 2367.100 210.000 ;
 END
END DIB83
PIN DOB83
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2352.960 208.880 2354.080 210.000 ;
  LAYER metal4 ;
  RECT 2352.960 208.880 2354.080 210.000 ;
  LAYER metal3 ;
  RECT 2352.960 208.880 2354.080 210.000 ;
  LAYER metal2 ;
  RECT 2352.960 208.880 2354.080 210.000 ;
  LAYER metal1 ;
  RECT 2352.960 208.880 2354.080 210.000 ;
 END
END DOB83
PIN DIB82
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2339.320 208.880 2340.440 210.000 ;
  LAYER metal4 ;
  RECT 2339.320 208.880 2340.440 210.000 ;
  LAYER metal3 ;
  RECT 2339.320 208.880 2340.440 210.000 ;
  LAYER metal2 ;
  RECT 2339.320 208.880 2340.440 210.000 ;
  LAYER metal1 ;
  RECT 2339.320 208.880 2340.440 210.000 ;
 END
END DIB82
PIN DOB82
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2325.680 208.880 2326.800 210.000 ;
  LAYER metal4 ;
  RECT 2325.680 208.880 2326.800 210.000 ;
  LAYER metal3 ;
  RECT 2325.680 208.880 2326.800 210.000 ;
  LAYER metal2 ;
  RECT 2325.680 208.880 2326.800 210.000 ;
  LAYER metal1 ;
  RECT 2325.680 208.880 2326.800 210.000 ;
 END
END DOB82
PIN DIB81
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2312.660 208.880 2313.780 210.000 ;
  LAYER metal4 ;
  RECT 2312.660 208.880 2313.780 210.000 ;
  LAYER metal3 ;
  RECT 2312.660 208.880 2313.780 210.000 ;
  LAYER metal2 ;
  RECT 2312.660 208.880 2313.780 210.000 ;
  LAYER metal1 ;
  RECT 2312.660 208.880 2313.780 210.000 ;
 END
END DIB81
PIN DOB81
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2299.020 208.880 2300.140 210.000 ;
  LAYER metal4 ;
  RECT 2299.020 208.880 2300.140 210.000 ;
  LAYER metal3 ;
  RECT 2299.020 208.880 2300.140 210.000 ;
  LAYER metal2 ;
  RECT 2299.020 208.880 2300.140 210.000 ;
  LAYER metal1 ;
  RECT 2299.020 208.880 2300.140 210.000 ;
 END
END DOB81
PIN DIB80
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2285.380 208.880 2286.500 210.000 ;
  LAYER metal4 ;
  RECT 2285.380 208.880 2286.500 210.000 ;
  LAYER metal3 ;
  RECT 2285.380 208.880 2286.500 210.000 ;
  LAYER metal2 ;
  RECT 2285.380 208.880 2286.500 210.000 ;
  LAYER metal1 ;
  RECT 2285.380 208.880 2286.500 210.000 ;
 END
END DIB80
PIN DOB80
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2272.360 208.880 2273.480 210.000 ;
  LAYER metal4 ;
  RECT 2272.360 208.880 2273.480 210.000 ;
  LAYER metal3 ;
  RECT 2272.360 208.880 2273.480 210.000 ;
  LAYER metal2 ;
  RECT 2272.360 208.880 2273.480 210.000 ;
  LAYER metal1 ;
  RECT 2272.360 208.880 2273.480 210.000 ;
 END
END DOB80
PIN DIB79
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2258.720 208.880 2259.840 210.000 ;
  LAYER metal4 ;
  RECT 2258.720 208.880 2259.840 210.000 ;
  LAYER metal3 ;
  RECT 2258.720 208.880 2259.840 210.000 ;
  LAYER metal2 ;
  RECT 2258.720 208.880 2259.840 210.000 ;
  LAYER metal1 ;
  RECT 2258.720 208.880 2259.840 210.000 ;
 END
END DIB79
PIN DOB79
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2245.080 208.880 2246.200 210.000 ;
  LAYER metal4 ;
  RECT 2245.080 208.880 2246.200 210.000 ;
  LAYER metal3 ;
  RECT 2245.080 208.880 2246.200 210.000 ;
  LAYER metal2 ;
  RECT 2245.080 208.880 2246.200 210.000 ;
  LAYER metal1 ;
  RECT 2245.080 208.880 2246.200 210.000 ;
 END
END DOB79
PIN DIB78
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2232.060 208.880 2233.180 210.000 ;
  LAYER metal4 ;
  RECT 2232.060 208.880 2233.180 210.000 ;
  LAYER metal3 ;
  RECT 2232.060 208.880 2233.180 210.000 ;
  LAYER metal2 ;
  RECT 2232.060 208.880 2233.180 210.000 ;
  LAYER metal1 ;
  RECT 2232.060 208.880 2233.180 210.000 ;
 END
END DIB78
PIN DOB78
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2218.420 208.880 2219.540 210.000 ;
  LAYER metal4 ;
  RECT 2218.420 208.880 2219.540 210.000 ;
  LAYER metal3 ;
  RECT 2218.420 208.880 2219.540 210.000 ;
  LAYER metal2 ;
  RECT 2218.420 208.880 2219.540 210.000 ;
  LAYER metal1 ;
  RECT 2218.420 208.880 2219.540 210.000 ;
 END
END DOB78
PIN DIB77
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2204.780 208.880 2205.900 210.000 ;
  LAYER metal4 ;
  RECT 2204.780 208.880 2205.900 210.000 ;
  LAYER metal3 ;
  RECT 2204.780 208.880 2205.900 210.000 ;
  LAYER metal2 ;
  RECT 2204.780 208.880 2205.900 210.000 ;
  LAYER metal1 ;
  RECT 2204.780 208.880 2205.900 210.000 ;
 END
END DIB77
PIN DOB77
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2191.140 208.880 2192.260 210.000 ;
  LAYER metal4 ;
  RECT 2191.140 208.880 2192.260 210.000 ;
  LAYER metal3 ;
  RECT 2191.140 208.880 2192.260 210.000 ;
  LAYER metal2 ;
  RECT 2191.140 208.880 2192.260 210.000 ;
  LAYER metal1 ;
  RECT 2191.140 208.880 2192.260 210.000 ;
 END
END DOB77
PIN DIB76
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2178.120 208.880 2179.240 210.000 ;
  LAYER metal4 ;
  RECT 2178.120 208.880 2179.240 210.000 ;
  LAYER metal3 ;
  RECT 2178.120 208.880 2179.240 210.000 ;
  LAYER metal2 ;
  RECT 2178.120 208.880 2179.240 210.000 ;
  LAYER metal1 ;
  RECT 2178.120 208.880 2179.240 210.000 ;
 END
END DIB76
PIN DOB76
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2164.480 208.880 2165.600 210.000 ;
  LAYER metal4 ;
  RECT 2164.480 208.880 2165.600 210.000 ;
  LAYER metal3 ;
  RECT 2164.480 208.880 2165.600 210.000 ;
  LAYER metal2 ;
  RECT 2164.480 208.880 2165.600 210.000 ;
  LAYER metal1 ;
  RECT 2164.480 208.880 2165.600 210.000 ;
 END
END DOB76
PIN DIB75
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2150.840 208.880 2151.960 210.000 ;
  LAYER metal4 ;
  RECT 2150.840 208.880 2151.960 210.000 ;
  LAYER metal3 ;
  RECT 2150.840 208.880 2151.960 210.000 ;
  LAYER metal2 ;
  RECT 2150.840 208.880 2151.960 210.000 ;
  LAYER metal1 ;
  RECT 2150.840 208.880 2151.960 210.000 ;
 END
END DIB75
PIN DOB75
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2137.820 208.880 2138.940 210.000 ;
  LAYER metal4 ;
  RECT 2137.820 208.880 2138.940 210.000 ;
  LAYER metal3 ;
  RECT 2137.820 208.880 2138.940 210.000 ;
  LAYER metal2 ;
  RECT 2137.820 208.880 2138.940 210.000 ;
  LAYER metal1 ;
  RECT 2137.820 208.880 2138.940 210.000 ;
 END
END DOB75
PIN DIB74
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2124.180 208.880 2125.300 210.000 ;
  LAYER metal4 ;
  RECT 2124.180 208.880 2125.300 210.000 ;
  LAYER metal3 ;
  RECT 2124.180 208.880 2125.300 210.000 ;
  LAYER metal2 ;
  RECT 2124.180 208.880 2125.300 210.000 ;
  LAYER metal1 ;
  RECT 2124.180 208.880 2125.300 210.000 ;
 END
END DIB74
PIN DOB74
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2110.540 208.880 2111.660 210.000 ;
  LAYER metal4 ;
  RECT 2110.540 208.880 2111.660 210.000 ;
  LAYER metal3 ;
  RECT 2110.540 208.880 2111.660 210.000 ;
  LAYER metal2 ;
  RECT 2110.540 208.880 2111.660 210.000 ;
  LAYER metal1 ;
  RECT 2110.540 208.880 2111.660 210.000 ;
 END
END DOB74
PIN DIB73
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2097.520 208.880 2098.640 210.000 ;
  LAYER metal4 ;
  RECT 2097.520 208.880 2098.640 210.000 ;
  LAYER metal3 ;
  RECT 2097.520 208.880 2098.640 210.000 ;
  LAYER metal2 ;
  RECT 2097.520 208.880 2098.640 210.000 ;
  LAYER metal1 ;
  RECT 2097.520 208.880 2098.640 210.000 ;
 END
END DIB73
PIN DOB73
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2083.880 208.880 2085.000 210.000 ;
  LAYER metal4 ;
  RECT 2083.880 208.880 2085.000 210.000 ;
  LAYER metal3 ;
  RECT 2083.880 208.880 2085.000 210.000 ;
  LAYER metal2 ;
  RECT 2083.880 208.880 2085.000 210.000 ;
  LAYER metal1 ;
  RECT 2083.880 208.880 2085.000 210.000 ;
 END
END DOB73
PIN DIB72
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2070.240 208.880 2071.360 210.000 ;
  LAYER metal4 ;
  RECT 2070.240 208.880 2071.360 210.000 ;
  LAYER metal3 ;
  RECT 2070.240 208.880 2071.360 210.000 ;
  LAYER metal2 ;
  RECT 2070.240 208.880 2071.360 210.000 ;
  LAYER metal1 ;
  RECT 2070.240 208.880 2071.360 210.000 ;
 END
END DIB72
PIN DOB72
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2057.220 208.880 2058.340 210.000 ;
  LAYER metal4 ;
  RECT 2057.220 208.880 2058.340 210.000 ;
  LAYER metal3 ;
  RECT 2057.220 208.880 2058.340 210.000 ;
  LAYER metal2 ;
  RECT 2057.220 208.880 2058.340 210.000 ;
  LAYER metal1 ;
  RECT 2057.220 208.880 2058.340 210.000 ;
 END
END DOB72
PIN DIB71
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2043.580 208.880 2044.700 210.000 ;
  LAYER metal4 ;
  RECT 2043.580 208.880 2044.700 210.000 ;
  LAYER metal3 ;
  RECT 2043.580 208.880 2044.700 210.000 ;
  LAYER metal2 ;
  RECT 2043.580 208.880 2044.700 210.000 ;
  LAYER metal1 ;
  RECT 2043.580 208.880 2044.700 210.000 ;
 END
END DIB71
PIN DOB71
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2029.940 208.880 2031.060 210.000 ;
  LAYER metal4 ;
  RECT 2029.940 208.880 2031.060 210.000 ;
  LAYER metal3 ;
  RECT 2029.940 208.880 2031.060 210.000 ;
  LAYER metal2 ;
  RECT 2029.940 208.880 2031.060 210.000 ;
  LAYER metal1 ;
  RECT 2029.940 208.880 2031.060 210.000 ;
 END
END DOB71
PIN DIB70
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2016.920 208.880 2018.040 210.000 ;
  LAYER metal4 ;
  RECT 2016.920 208.880 2018.040 210.000 ;
  LAYER metal3 ;
  RECT 2016.920 208.880 2018.040 210.000 ;
  LAYER metal2 ;
  RECT 2016.920 208.880 2018.040 210.000 ;
  LAYER metal1 ;
  RECT 2016.920 208.880 2018.040 210.000 ;
 END
END DIB70
PIN DOB70
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2003.280 208.880 2004.400 210.000 ;
  LAYER metal4 ;
  RECT 2003.280 208.880 2004.400 210.000 ;
  LAYER metal3 ;
  RECT 2003.280 208.880 2004.400 210.000 ;
  LAYER metal2 ;
  RECT 2003.280 208.880 2004.400 210.000 ;
  LAYER metal1 ;
  RECT 2003.280 208.880 2004.400 210.000 ;
 END
END DOB70
PIN DIB69
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1989.640 208.880 1990.760 210.000 ;
  LAYER metal4 ;
  RECT 1989.640 208.880 1990.760 210.000 ;
  LAYER metal3 ;
  RECT 1989.640 208.880 1990.760 210.000 ;
  LAYER metal2 ;
  RECT 1989.640 208.880 1990.760 210.000 ;
  LAYER metal1 ;
  RECT 1989.640 208.880 1990.760 210.000 ;
 END
END DIB69
PIN DOB69
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1976.620 208.880 1977.740 210.000 ;
  LAYER metal4 ;
  RECT 1976.620 208.880 1977.740 210.000 ;
  LAYER metal3 ;
  RECT 1976.620 208.880 1977.740 210.000 ;
  LAYER metal2 ;
  RECT 1976.620 208.880 1977.740 210.000 ;
  LAYER metal1 ;
  RECT 1976.620 208.880 1977.740 210.000 ;
 END
END DOB69
PIN DIB68
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1962.980 208.880 1964.100 210.000 ;
  LAYER metal4 ;
  RECT 1962.980 208.880 1964.100 210.000 ;
  LAYER metal3 ;
  RECT 1962.980 208.880 1964.100 210.000 ;
  LAYER metal2 ;
  RECT 1962.980 208.880 1964.100 210.000 ;
  LAYER metal1 ;
  RECT 1962.980 208.880 1964.100 210.000 ;
 END
END DIB68
PIN DOB68
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1949.340 208.880 1950.460 210.000 ;
  LAYER metal4 ;
  RECT 1949.340 208.880 1950.460 210.000 ;
  LAYER metal3 ;
  RECT 1949.340 208.880 1950.460 210.000 ;
  LAYER metal2 ;
  RECT 1949.340 208.880 1950.460 210.000 ;
  LAYER metal1 ;
  RECT 1949.340 208.880 1950.460 210.000 ;
 END
END DOB68
PIN DIB67
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1936.320 208.880 1937.440 210.000 ;
  LAYER metal4 ;
  RECT 1936.320 208.880 1937.440 210.000 ;
  LAYER metal3 ;
  RECT 1936.320 208.880 1937.440 210.000 ;
  LAYER metal2 ;
  RECT 1936.320 208.880 1937.440 210.000 ;
  LAYER metal1 ;
  RECT 1936.320 208.880 1937.440 210.000 ;
 END
END DIB67
PIN DOB67
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1922.680 208.880 1923.800 210.000 ;
  LAYER metal4 ;
  RECT 1922.680 208.880 1923.800 210.000 ;
  LAYER metal3 ;
  RECT 1922.680 208.880 1923.800 210.000 ;
  LAYER metal2 ;
  RECT 1922.680 208.880 1923.800 210.000 ;
  LAYER metal1 ;
  RECT 1922.680 208.880 1923.800 210.000 ;
 END
END DOB67
PIN DIB66
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1909.040 208.880 1910.160 210.000 ;
  LAYER metal4 ;
  RECT 1909.040 208.880 1910.160 210.000 ;
  LAYER metal3 ;
  RECT 1909.040 208.880 1910.160 210.000 ;
  LAYER metal2 ;
  RECT 1909.040 208.880 1910.160 210.000 ;
  LAYER metal1 ;
  RECT 1909.040 208.880 1910.160 210.000 ;
 END
END DIB66
PIN DOB66
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1896.020 208.880 1897.140 210.000 ;
  LAYER metal4 ;
  RECT 1896.020 208.880 1897.140 210.000 ;
  LAYER metal3 ;
  RECT 1896.020 208.880 1897.140 210.000 ;
  LAYER metal2 ;
  RECT 1896.020 208.880 1897.140 210.000 ;
  LAYER metal1 ;
  RECT 1896.020 208.880 1897.140 210.000 ;
 END
END DOB66
PIN DIB65
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1882.380 208.880 1883.500 210.000 ;
  LAYER metal4 ;
  RECT 1882.380 208.880 1883.500 210.000 ;
  LAYER metal3 ;
  RECT 1882.380 208.880 1883.500 210.000 ;
  LAYER metal2 ;
  RECT 1882.380 208.880 1883.500 210.000 ;
  LAYER metal1 ;
  RECT 1882.380 208.880 1883.500 210.000 ;
 END
END DIB65
PIN DOB65
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1868.740 208.880 1869.860 210.000 ;
  LAYER metal4 ;
  RECT 1868.740 208.880 1869.860 210.000 ;
  LAYER metal3 ;
  RECT 1868.740 208.880 1869.860 210.000 ;
  LAYER metal2 ;
  RECT 1868.740 208.880 1869.860 210.000 ;
  LAYER metal1 ;
  RECT 1868.740 208.880 1869.860 210.000 ;
 END
END DOB65
PIN DIB64
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1855.720 208.880 1856.840 210.000 ;
  LAYER metal4 ;
  RECT 1855.720 208.880 1856.840 210.000 ;
  LAYER metal3 ;
  RECT 1855.720 208.880 1856.840 210.000 ;
  LAYER metal2 ;
  RECT 1855.720 208.880 1856.840 210.000 ;
  LAYER metal1 ;
  RECT 1855.720 208.880 1856.840 210.000 ;
 END
END DIB64
PIN DOB64
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1842.080 208.880 1843.200 210.000 ;
  LAYER metal4 ;
  RECT 1842.080 208.880 1843.200 210.000 ;
  LAYER metal3 ;
  RECT 1842.080 208.880 1843.200 210.000 ;
  LAYER metal2 ;
  RECT 1842.080 208.880 1843.200 210.000 ;
  LAYER metal1 ;
  RECT 1842.080 208.880 1843.200 210.000 ;
 END
END DOB64
PIN OEB
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1815.420 208.880 1816.540 210.000 ;
  LAYER metal4 ;
  RECT 1815.420 208.880 1816.540 210.000 ;
  LAYER metal3 ;
  RECT 1815.420 208.880 1816.540 210.000 ;
  LAYER metal2 ;
  RECT 1815.420 208.880 1816.540 210.000 ;
  LAYER metal1 ;
  RECT 1815.420 208.880 1816.540 210.000 ;
 END
END OEB
PIN CKB
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1801.780 208.880 1802.900 210.000 ;
  LAYER metal4 ;
  RECT 1801.780 208.880 1802.900 210.000 ;
  LAYER metal3 ;
  RECT 1801.780 208.880 1802.900 210.000 ;
  LAYER metal2 ;
  RECT 1801.780 208.880 1802.900 210.000 ;
  LAYER metal1 ;
  RECT 1801.780 208.880 1802.900 210.000 ;
 END
END CKB
PIN CSB
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1799.920 208.880 1801.040 210.000 ;
  LAYER metal4 ;
  RECT 1799.920 208.880 1801.040 210.000 ;
  LAYER metal3 ;
  RECT 1799.920 208.880 1801.040 210.000 ;
  LAYER metal2 ;
  RECT 1799.920 208.880 1801.040 210.000 ;
  LAYER metal1 ;
  RECT 1799.920 208.880 1801.040 210.000 ;
 END
END CSB
PIN WEBN
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1797.440 208.880 1798.560 210.000 ;
  LAYER metal4 ;
  RECT 1797.440 208.880 1798.560 210.000 ;
  LAYER metal3 ;
  RECT 1797.440 208.880 1798.560 210.000 ;
  LAYER metal2 ;
  RECT 1797.440 208.880 1798.560 210.000 ;
  LAYER metal1 ;
  RECT 1797.440 208.880 1798.560 210.000 ;
 END
END WEBN
PIN B2
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1793.720 208.880 1794.840 210.000 ;
  LAYER metal4 ;
  RECT 1793.720 208.880 1794.840 210.000 ;
  LAYER metal3 ;
  RECT 1793.720 208.880 1794.840 210.000 ;
  LAYER metal2 ;
  RECT 1793.720 208.880 1794.840 210.000 ;
  LAYER metal1 ;
  RECT 1793.720 208.880 1794.840 210.000 ;
 END
END B2
PIN B1
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1788.140 208.880 1789.260 210.000 ;
  LAYER metal4 ;
  RECT 1788.140 208.880 1789.260 210.000 ;
  LAYER metal3 ;
  RECT 1788.140 208.880 1789.260 210.000 ;
  LAYER metal2 ;
  RECT 1788.140 208.880 1789.260 210.000 ;
  LAYER metal1 ;
  RECT 1788.140 208.880 1789.260 210.000 ;
 END
END B1
PIN B0
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1786.280 208.880 1787.400 210.000 ;
  LAYER metal4 ;
  RECT 1786.280 208.880 1787.400 210.000 ;
  LAYER metal3 ;
  RECT 1786.280 208.880 1787.400 210.000 ;
  LAYER metal2 ;
  RECT 1786.280 208.880 1787.400 210.000 ;
  LAYER metal1 ;
  RECT 1786.280 208.880 1787.400 210.000 ;
 END
END B0
PIN B5
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1777.600 208.880 1778.720 210.000 ;
  LAYER metal4 ;
  RECT 1777.600 208.880 1778.720 210.000 ;
  LAYER metal3 ;
  RECT 1777.600 208.880 1778.720 210.000 ;
  LAYER metal2 ;
  RECT 1777.600 208.880 1778.720 210.000 ;
  LAYER metal1 ;
  RECT 1777.600 208.880 1778.720 210.000 ;
 END
END B5
PIN B4
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1772.020 208.880 1773.140 210.000 ;
  LAYER metal4 ;
  RECT 1772.020 208.880 1773.140 210.000 ;
  LAYER metal3 ;
  RECT 1772.020 208.880 1773.140 210.000 ;
  LAYER metal2 ;
  RECT 1772.020 208.880 1773.140 210.000 ;
  LAYER metal1 ;
  RECT 1772.020 208.880 1773.140 210.000 ;
 END
END B4
PIN B3
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1766.440 208.880 1767.560 210.000 ;
  LAYER metal4 ;
  RECT 1766.440 208.880 1767.560 210.000 ;
  LAYER metal3 ;
  RECT 1766.440 208.880 1767.560 210.000 ;
  LAYER metal2 ;
  RECT 1766.440 208.880 1767.560 210.000 ;
  LAYER metal1 ;
  RECT 1766.440 208.880 1767.560 210.000 ;
 END
END B3
PIN B7
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1747.840 208.880 1748.960 210.000 ;
  LAYER metal4 ;
  RECT 1747.840 208.880 1748.960 210.000 ;
  LAYER metal3 ;
  RECT 1747.840 208.880 1748.960 210.000 ;
  LAYER metal2 ;
  RECT 1747.840 208.880 1748.960 210.000 ;
  LAYER metal1 ;
  RECT 1747.840 208.880 1748.960 210.000 ;
 END
END B7
PIN B6
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1741.640 208.880 1742.760 210.000 ;
  LAYER metal4 ;
  RECT 1741.640 208.880 1742.760 210.000 ;
  LAYER metal3 ;
  RECT 1741.640 208.880 1742.760 210.000 ;
  LAYER metal2 ;
  RECT 1741.640 208.880 1742.760 210.000 ;
  LAYER metal1 ;
  RECT 1741.640 208.880 1742.760 210.000 ;
 END
END B6
PIN DIB63
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1719.320 208.880 1720.440 210.000 ;
  LAYER metal4 ;
  RECT 1719.320 208.880 1720.440 210.000 ;
  LAYER metal3 ;
  RECT 1719.320 208.880 1720.440 210.000 ;
  LAYER metal2 ;
  RECT 1719.320 208.880 1720.440 210.000 ;
  LAYER metal1 ;
  RECT 1719.320 208.880 1720.440 210.000 ;
 END
END DIB63
PIN DOB63
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1706.300 208.880 1707.420 210.000 ;
  LAYER metal4 ;
  RECT 1706.300 208.880 1707.420 210.000 ;
  LAYER metal3 ;
  RECT 1706.300 208.880 1707.420 210.000 ;
  LAYER metal2 ;
  RECT 1706.300 208.880 1707.420 210.000 ;
  LAYER metal1 ;
  RECT 1706.300 208.880 1707.420 210.000 ;
 END
END DOB63
PIN DIB62
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1692.660 208.880 1693.780 210.000 ;
  LAYER metal4 ;
  RECT 1692.660 208.880 1693.780 210.000 ;
  LAYER metal3 ;
  RECT 1692.660 208.880 1693.780 210.000 ;
  LAYER metal2 ;
  RECT 1692.660 208.880 1693.780 210.000 ;
  LAYER metal1 ;
  RECT 1692.660 208.880 1693.780 210.000 ;
 END
END DIB62
PIN DOB62
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1679.020 208.880 1680.140 210.000 ;
  LAYER metal4 ;
  RECT 1679.020 208.880 1680.140 210.000 ;
  LAYER metal3 ;
  RECT 1679.020 208.880 1680.140 210.000 ;
  LAYER metal2 ;
  RECT 1679.020 208.880 1680.140 210.000 ;
  LAYER metal1 ;
  RECT 1679.020 208.880 1680.140 210.000 ;
 END
END DOB62
PIN DIB61
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1666.000 208.880 1667.120 210.000 ;
  LAYER metal4 ;
  RECT 1666.000 208.880 1667.120 210.000 ;
  LAYER metal3 ;
  RECT 1666.000 208.880 1667.120 210.000 ;
  LAYER metal2 ;
  RECT 1666.000 208.880 1667.120 210.000 ;
  LAYER metal1 ;
  RECT 1666.000 208.880 1667.120 210.000 ;
 END
END DIB61
PIN DOB61
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1652.360 208.880 1653.480 210.000 ;
  LAYER metal4 ;
  RECT 1652.360 208.880 1653.480 210.000 ;
  LAYER metal3 ;
  RECT 1652.360 208.880 1653.480 210.000 ;
  LAYER metal2 ;
  RECT 1652.360 208.880 1653.480 210.000 ;
  LAYER metal1 ;
  RECT 1652.360 208.880 1653.480 210.000 ;
 END
END DOB61
PIN DIB60
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1638.720 208.880 1639.840 210.000 ;
  LAYER metal4 ;
  RECT 1638.720 208.880 1639.840 210.000 ;
  LAYER metal3 ;
  RECT 1638.720 208.880 1639.840 210.000 ;
  LAYER metal2 ;
  RECT 1638.720 208.880 1639.840 210.000 ;
  LAYER metal1 ;
  RECT 1638.720 208.880 1639.840 210.000 ;
 END
END DIB60
PIN DOB60
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1625.700 208.880 1626.820 210.000 ;
  LAYER metal4 ;
  RECT 1625.700 208.880 1626.820 210.000 ;
  LAYER metal3 ;
  RECT 1625.700 208.880 1626.820 210.000 ;
  LAYER metal2 ;
  RECT 1625.700 208.880 1626.820 210.000 ;
  LAYER metal1 ;
  RECT 1625.700 208.880 1626.820 210.000 ;
 END
END DOB60
PIN DIB59
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1612.060 208.880 1613.180 210.000 ;
  LAYER metal4 ;
  RECT 1612.060 208.880 1613.180 210.000 ;
  LAYER metal3 ;
  RECT 1612.060 208.880 1613.180 210.000 ;
  LAYER metal2 ;
  RECT 1612.060 208.880 1613.180 210.000 ;
  LAYER metal1 ;
  RECT 1612.060 208.880 1613.180 210.000 ;
 END
END DIB59
PIN DOB59
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1598.420 208.880 1599.540 210.000 ;
  LAYER metal4 ;
  RECT 1598.420 208.880 1599.540 210.000 ;
  LAYER metal3 ;
  RECT 1598.420 208.880 1599.540 210.000 ;
  LAYER metal2 ;
  RECT 1598.420 208.880 1599.540 210.000 ;
  LAYER metal1 ;
  RECT 1598.420 208.880 1599.540 210.000 ;
 END
END DOB59
PIN DIB58
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1585.400 208.880 1586.520 210.000 ;
  LAYER metal4 ;
  RECT 1585.400 208.880 1586.520 210.000 ;
  LAYER metal3 ;
  RECT 1585.400 208.880 1586.520 210.000 ;
  LAYER metal2 ;
  RECT 1585.400 208.880 1586.520 210.000 ;
  LAYER metal1 ;
  RECT 1585.400 208.880 1586.520 210.000 ;
 END
END DIB58
PIN DOB58
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1571.760 208.880 1572.880 210.000 ;
  LAYER metal4 ;
  RECT 1571.760 208.880 1572.880 210.000 ;
  LAYER metal3 ;
  RECT 1571.760 208.880 1572.880 210.000 ;
  LAYER metal2 ;
  RECT 1571.760 208.880 1572.880 210.000 ;
  LAYER metal1 ;
  RECT 1571.760 208.880 1572.880 210.000 ;
 END
END DOB58
PIN DIB57
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1558.120 208.880 1559.240 210.000 ;
  LAYER metal4 ;
  RECT 1558.120 208.880 1559.240 210.000 ;
  LAYER metal3 ;
  RECT 1558.120 208.880 1559.240 210.000 ;
  LAYER metal2 ;
  RECT 1558.120 208.880 1559.240 210.000 ;
  LAYER metal1 ;
  RECT 1558.120 208.880 1559.240 210.000 ;
 END
END DIB57
PIN DOB57
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1545.100 208.880 1546.220 210.000 ;
  LAYER metal4 ;
  RECT 1545.100 208.880 1546.220 210.000 ;
  LAYER metal3 ;
  RECT 1545.100 208.880 1546.220 210.000 ;
  LAYER metal2 ;
  RECT 1545.100 208.880 1546.220 210.000 ;
  LAYER metal1 ;
  RECT 1545.100 208.880 1546.220 210.000 ;
 END
END DOB57
PIN DIB56
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1531.460 208.880 1532.580 210.000 ;
  LAYER metal4 ;
  RECT 1531.460 208.880 1532.580 210.000 ;
  LAYER metal3 ;
  RECT 1531.460 208.880 1532.580 210.000 ;
  LAYER metal2 ;
  RECT 1531.460 208.880 1532.580 210.000 ;
  LAYER metal1 ;
  RECT 1531.460 208.880 1532.580 210.000 ;
 END
END DIB56
PIN DOB56
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1517.820 208.880 1518.940 210.000 ;
  LAYER metal4 ;
  RECT 1517.820 208.880 1518.940 210.000 ;
  LAYER metal3 ;
  RECT 1517.820 208.880 1518.940 210.000 ;
  LAYER metal2 ;
  RECT 1517.820 208.880 1518.940 210.000 ;
  LAYER metal1 ;
  RECT 1517.820 208.880 1518.940 210.000 ;
 END
END DOB56
PIN DIB55
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1504.800 208.880 1505.920 210.000 ;
  LAYER metal4 ;
  RECT 1504.800 208.880 1505.920 210.000 ;
  LAYER metal3 ;
  RECT 1504.800 208.880 1505.920 210.000 ;
  LAYER metal2 ;
  RECT 1504.800 208.880 1505.920 210.000 ;
  LAYER metal1 ;
  RECT 1504.800 208.880 1505.920 210.000 ;
 END
END DIB55
PIN DOB55
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1491.160 208.880 1492.280 210.000 ;
  LAYER metal4 ;
  RECT 1491.160 208.880 1492.280 210.000 ;
  LAYER metal3 ;
  RECT 1491.160 208.880 1492.280 210.000 ;
  LAYER metal2 ;
  RECT 1491.160 208.880 1492.280 210.000 ;
  LAYER metal1 ;
  RECT 1491.160 208.880 1492.280 210.000 ;
 END
END DOB55
PIN DIB54
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1477.520 208.880 1478.640 210.000 ;
  LAYER metal4 ;
  RECT 1477.520 208.880 1478.640 210.000 ;
  LAYER metal3 ;
  RECT 1477.520 208.880 1478.640 210.000 ;
  LAYER metal2 ;
  RECT 1477.520 208.880 1478.640 210.000 ;
  LAYER metal1 ;
  RECT 1477.520 208.880 1478.640 210.000 ;
 END
END DIB54
PIN DOB54
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1464.500 208.880 1465.620 210.000 ;
  LAYER metal4 ;
  RECT 1464.500 208.880 1465.620 210.000 ;
  LAYER metal3 ;
  RECT 1464.500 208.880 1465.620 210.000 ;
  LAYER metal2 ;
  RECT 1464.500 208.880 1465.620 210.000 ;
  LAYER metal1 ;
  RECT 1464.500 208.880 1465.620 210.000 ;
 END
END DOB54
PIN DIB53
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1450.860 208.880 1451.980 210.000 ;
  LAYER metal4 ;
  RECT 1450.860 208.880 1451.980 210.000 ;
  LAYER metal3 ;
  RECT 1450.860 208.880 1451.980 210.000 ;
  LAYER metal2 ;
  RECT 1450.860 208.880 1451.980 210.000 ;
  LAYER metal1 ;
  RECT 1450.860 208.880 1451.980 210.000 ;
 END
END DIB53
PIN DOB53
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1437.220 208.880 1438.340 210.000 ;
  LAYER metal4 ;
  RECT 1437.220 208.880 1438.340 210.000 ;
  LAYER metal3 ;
  RECT 1437.220 208.880 1438.340 210.000 ;
  LAYER metal2 ;
  RECT 1437.220 208.880 1438.340 210.000 ;
  LAYER metal1 ;
  RECT 1437.220 208.880 1438.340 210.000 ;
 END
END DOB53
PIN DIB52
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1424.200 208.880 1425.320 210.000 ;
  LAYER metal4 ;
  RECT 1424.200 208.880 1425.320 210.000 ;
  LAYER metal3 ;
  RECT 1424.200 208.880 1425.320 210.000 ;
  LAYER metal2 ;
  RECT 1424.200 208.880 1425.320 210.000 ;
  LAYER metal1 ;
  RECT 1424.200 208.880 1425.320 210.000 ;
 END
END DIB52
PIN DOB52
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1410.560 208.880 1411.680 210.000 ;
  LAYER metal4 ;
  RECT 1410.560 208.880 1411.680 210.000 ;
  LAYER metal3 ;
  RECT 1410.560 208.880 1411.680 210.000 ;
  LAYER metal2 ;
  RECT 1410.560 208.880 1411.680 210.000 ;
  LAYER metal1 ;
  RECT 1410.560 208.880 1411.680 210.000 ;
 END
END DOB52
PIN DIB51
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1396.920 208.880 1398.040 210.000 ;
  LAYER metal4 ;
  RECT 1396.920 208.880 1398.040 210.000 ;
  LAYER metal3 ;
  RECT 1396.920 208.880 1398.040 210.000 ;
  LAYER metal2 ;
  RECT 1396.920 208.880 1398.040 210.000 ;
  LAYER metal1 ;
  RECT 1396.920 208.880 1398.040 210.000 ;
 END
END DIB51
PIN DOB51
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1383.900 208.880 1385.020 210.000 ;
  LAYER metal4 ;
  RECT 1383.900 208.880 1385.020 210.000 ;
  LAYER metal3 ;
  RECT 1383.900 208.880 1385.020 210.000 ;
  LAYER metal2 ;
  RECT 1383.900 208.880 1385.020 210.000 ;
  LAYER metal1 ;
  RECT 1383.900 208.880 1385.020 210.000 ;
 END
END DOB51
PIN DIB50
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1370.260 208.880 1371.380 210.000 ;
  LAYER metal4 ;
  RECT 1370.260 208.880 1371.380 210.000 ;
  LAYER metal3 ;
  RECT 1370.260 208.880 1371.380 210.000 ;
  LAYER metal2 ;
  RECT 1370.260 208.880 1371.380 210.000 ;
  LAYER metal1 ;
  RECT 1370.260 208.880 1371.380 210.000 ;
 END
END DIB50
PIN DOB50
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1356.620 208.880 1357.740 210.000 ;
  LAYER metal4 ;
  RECT 1356.620 208.880 1357.740 210.000 ;
  LAYER metal3 ;
  RECT 1356.620 208.880 1357.740 210.000 ;
  LAYER metal2 ;
  RECT 1356.620 208.880 1357.740 210.000 ;
  LAYER metal1 ;
  RECT 1356.620 208.880 1357.740 210.000 ;
 END
END DOB50
PIN DIB49
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1343.600 208.880 1344.720 210.000 ;
  LAYER metal4 ;
  RECT 1343.600 208.880 1344.720 210.000 ;
  LAYER metal3 ;
  RECT 1343.600 208.880 1344.720 210.000 ;
  LAYER metal2 ;
  RECT 1343.600 208.880 1344.720 210.000 ;
  LAYER metal1 ;
  RECT 1343.600 208.880 1344.720 210.000 ;
 END
END DIB49
PIN DOB49
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1329.960 208.880 1331.080 210.000 ;
  LAYER metal4 ;
  RECT 1329.960 208.880 1331.080 210.000 ;
  LAYER metal3 ;
  RECT 1329.960 208.880 1331.080 210.000 ;
  LAYER metal2 ;
  RECT 1329.960 208.880 1331.080 210.000 ;
  LAYER metal1 ;
  RECT 1329.960 208.880 1331.080 210.000 ;
 END
END DOB49
PIN DIB48
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1316.320 208.880 1317.440 210.000 ;
  LAYER metal4 ;
  RECT 1316.320 208.880 1317.440 210.000 ;
  LAYER metal3 ;
  RECT 1316.320 208.880 1317.440 210.000 ;
  LAYER metal2 ;
  RECT 1316.320 208.880 1317.440 210.000 ;
  LAYER metal1 ;
  RECT 1316.320 208.880 1317.440 210.000 ;
 END
END DIB48
PIN DOB48
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1302.680 208.880 1303.800 210.000 ;
  LAYER metal4 ;
  RECT 1302.680 208.880 1303.800 210.000 ;
  LAYER metal3 ;
  RECT 1302.680 208.880 1303.800 210.000 ;
  LAYER metal2 ;
  RECT 1302.680 208.880 1303.800 210.000 ;
  LAYER metal1 ;
  RECT 1302.680 208.880 1303.800 210.000 ;
 END
END DOB48
PIN DIB47
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1289.660 208.880 1290.780 210.000 ;
  LAYER metal4 ;
  RECT 1289.660 208.880 1290.780 210.000 ;
  LAYER metal3 ;
  RECT 1289.660 208.880 1290.780 210.000 ;
  LAYER metal2 ;
  RECT 1289.660 208.880 1290.780 210.000 ;
  LAYER metal1 ;
  RECT 1289.660 208.880 1290.780 210.000 ;
 END
END DIB47
PIN DOB47
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1276.020 208.880 1277.140 210.000 ;
  LAYER metal4 ;
  RECT 1276.020 208.880 1277.140 210.000 ;
  LAYER metal3 ;
  RECT 1276.020 208.880 1277.140 210.000 ;
  LAYER metal2 ;
  RECT 1276.020 208.880 1277.140 210.000 ;
  LAYER metal1 ;
  RECT 1276.020 208.880 1277.140 210.000 ;
 END
END DOB47
PIN DIB46
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1262.380 208.880 1263.500 210.000 ;
  LAYER metal4 ;
  RECT 1262.380 208.880 1263.500 210.000 ;
  LAYER metal3 ;
  RECT 1262.380 208.880 1263.500 210.000 ;
  LAYER metal2 ;
  RECT 1262.380 208.880 1263.500 210.000 ;
  LAYER metal1 ;
  RECT 1262.380 208.880 1263.500 210.000 ;
 END
END DIB46
PIN DOB46
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1249.360 208.880 1250.480 210.000 ;
  LAYER metal4 ;
  RECT 1249.360 208.880 1250.480 210.000 ;
  LAYER metal3 ;
  RECT 1249.360 208.880 1250.480 210.000 ;
  LAYER metal2 ;
  RECT 1249.360 208.880 1250.480 210.000 ;
  LAYER metal1 ;
  RECT 1249.360 208.880 1250.480 210.000 ;
 END
END DOB46
PIN DIB45
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1235.720 208.880 1236.840 210.000 ;
  LAYER metal4 ;
  RECT 1235.720 208.880 1236.840 210.000 ;
  LAYER metal3 ;
  RECT 1235.720 208.880 1236.840 210.000 ;
  LAYER metal2 ;
  RECT 1235.720 208.880 1236.840 210.000 ;
  LAYER metal1 ;
  RECT 1235.720 208.880 1236.840 210.000 ;
 END
END DIB45
PIN DOB45
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1222.080 208.880 1223.200 210.000 ;
  LAYER metal4 ;
  RECT 1222.080 208.880 1223.200 210.000 ;
  LAYER metal3 ;
  RECT 1222.080 208.880 1223.200 210.000 ;
  LAYER metal2 ;
  RECT 1222.080 208.880 1223.200 210.000 ;
  LAYER metal1 ;
  RECT 1222.080 208.880 1223.200 210.000 ;
 END
END DOB45
PIN DIB44
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1209.060 208.880 1210.180 210.000 ;
  LAYER metal4 ;
  RECT 1209.060 208.880 1210.180 210.000 ;
  LAYER metal3 ;
  RECT 1209.060 208.880 1210.180 210.000 ;
  LAYER metal2 ;
  RECT 1209.060 208.880 1210.180 210.000 ;
  LAYER metal1 ;
  RECT 1209.060 208.880 1210.180 210.000 ;
 END
END DIB44
PIN DOB44
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1195.420 208.880 1196.540 210.000 ;
  LAYER metal4 ;
  RECT 1195.420 208.880 1196.540 210.000 ;
  LAYER metal3 ;
  RECT 1195.420 208.880 1196.540 210.000 ;
  LAYER metal2 ;
  RECT 1195.420 208.880 1196.540 210.000 ;
  LAYER metal1 ;
  RECT 1195.420 208.880 1196.540 210.000 ;
 END
END DOB44
PIN DIB43
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1181.780 208.880 1182.900 210.000 ;
  LAYER metal4 ;
  RECT 1181.780 208.880 1182.900 210.000 ;
  LAYER metal3 ;
  RECT 1181.780 208.880 1182.900 210.000 ;
  LAYER metal2 ;
  RECT 1181.780 208.880 1182.900 210.000 ;
  LAYER metal1 ;
  RECT 1181.780 208.880 1182.900 210.000 ;
 END
END DIB43
PIN DOB43
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1168.760 208.880 1169.880 210.000 ;
  LAYER metal4 ;
  RECT 1168.760 208.880 1169.880 210.000 ;
  LAYER metal3 ;
  RECT 1168.760 208.880 1169.880 210.000 ;
  LAYER metal2 ;
  RECT 1168.760 208.880 1169.880 210.000 ;
  LAYER metal1 ;
  RECT 1168.760 208.880 1169.880 210.000 ;
 END
END DOB43
PIN DIB42
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1155.120 208.880 1156.240 210.000 ;
  LAYER metal4 ;
  RECT 1155.120 208.880 1156.240 210.000 ;
  LAYER metal3 ;
  RECT 1155.120 208.880 1156.240 210.000 ;
  LAYER metal2 ;
  RECT 1155.120 208.880 1156.240 210.000 ;
  LAYER metal1 ;
  RECT 1155.120 208.880 1156.240 210.000 ;
 END
END DIB42
PIN DOB42
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1141.480 208.880 1142.600 210.000 ;
  LAYER metal4 ;
  RECT 1141.480 208.880 1142.600 210.000 ;
  LAYER metal3 ;
  RECT 1141.480 208.880 1142.600 210.000 ;
  LAYER metal2 ;
  RECT 1141.480 208.880 1142.600 210.000 ;
  LAYER metal1 ;
  RECT 1141.480 208.880 1142.600 210.000 ;
 END
END DOB42
PIN DIB41
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1128.460 208.880 1129.580 210.000 ;
  LAYER metal4 ;
  RECT 1128.460 208.880 1129.580 210.000 ;
  LAYER metal3 ;
  RECT 1128.460 208.880 1129.580 210.000 ;
  LAYER metal2 ;
  RECT 1128.460 208.880 1129.580 210.000 ;
  LAYER metal1 ;
  RECT 1128.460 208.880 1129.580 210.000 ;
 END
END DIB41
PIN DOB41
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1114.820 208.880 1115.940 210.000 ;
  LAYER metal4 ;
  RECT 1114.820 208.880 1115.940 210.000 ;
  LAYER metal3 ;
  RECT 1114.820 208.880 1115.940 210.000 ;
  LAYER metal2 ;
  RECT 1114.820 208.880 1115.940 210.000 ;
  LAYER metal1 ;
  RECT 1114.820 208.880 1115.940 210.000 ;
 END
END DOB41
PIN DIB40
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1101.180 208.880 1102.300 210.000 ;
  LAYER metal4 ;
  RECT 1101.180 208.880 1102.300 210.000 ;
  LAYER metal3 ;
  RECT 1101.180 208.880 1102.300 210.000 ;
  LAYER metal2 ;
  RECT 1101.180 208.880 1102.300 210.000 ;
  LAYER metal1 ;
  RECT 1101.180 208.880 1102.300 210.000 ;
 END
END DIB40
PIN DOB40
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1088.160 208.880 1089.280 210.000 ;
  LAYER metal4 ;
  RECT 1088.160 208.880 1089.280 210.000 ;
  LAYER metal3 ;
  RECT 1088.160 208.880 1089.280 210.000 ;
  LAYER metal2 ;
  RECT 1088.160 208.880 1089.280 210.000 ;
  LAYER metal1 ;
  RECT 1088.160 208.880 1089.280 210.000 ;
 END
END DOB40
PIN DIB39
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1074.520 208.880 1075.640 210.000 ;
  LAYER metal4 ;
  RECT 1074.520 208.880 1075.640 210.000 ;
  LAYER metal3 ;
  RECT 1074.520 208.880 1075.640 210.000 ;
  LAYER metal2 ;
  RECT 1074.520 208.880 1075.640 210.000 ;
  LAYER metal1 ;
  RECT 1074.520 208.880 1075.640 210.000 ;
 END
END DIB39
PIN DOB39
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1060.880 208.880 1062.000 210.000 ;
  LAYER metal4 ;
  RECT 1060.880 208.880 1062.000 210.000 ;
  LAYER metal3 ;
  RECT 1060.880 208.880 1062.000 210.000 ;
  LAYER metal2 ;
  RECT 1060.880 208.880 1062.000 210.000 ;
  LAYER metal1 ;
  RECT 1060.880 208.880 1062.000 210.000 ;
 END
END DOB39
PIN DIB38
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1047.860 208.880 1048.980 210.000 ;
  LAYER metal4 ;
  RECT 1047.860 208.880 1048.980 210.000 ;
  LAYER metal3 ;
  RECT 1047.860 208.880 1048.980 210.000 ;
  LAYER metal2 ;
  RECT 1047.860 208.880 1048.980 210.000 ;
  LAYER metal1 ;
  RECT 1047.860 208.880 1048.980 210.000 ;
 END
END DIB38
PIN DOB38
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1034.220 208.880 1035.340 210.000 ;
  LAYER metal4 ;
  RECT 1034.220 208.880 1035.340 210.000 ;
  LAYER metal3 ;
  RECT 1034.220 208.880 1035.340 210.000 ;
  LAYER metal2 ;
  RECT 1034.220 208.880 1035.340 210.000 ;
  LAYER metal1 ;
  RECT 1034.220 208.880 1035.340 210.000 ;
 END
END DOB38
PIN DIB37
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1020.580 208.880 1021.700 210.000 ;
  LAYER metal4 ;
  RECT 1020.580 208.880 1021.700 210.000 ;
  LAYER metal3 ;
  RECT 1020.580 208.880 1021.700 210.000 ;
  LAYER metal2 ;
  RECT 1020.580 208.880 1021.700 210.000 ;
  LAYER metal1 ;
  RECT 1020.580 208.880 1021.700 210.000 ;
 END
END DIB37
PIN DOB37
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1007.560 208.880 1008.680 210.000 ;
  LAYER metal4 ;
  RECT 1007.560 208.880 1008.680 210.000 ;
  LAYER metal3 ;
  RECT 1007.560 208.880 1008.680 210.000 ;
  LAYER metal2 ;
  RECT 1007.560 208.880 1008.680 210.000 ;
  LAYER metal1 ;
  RECT 1007.560 208.880 1008.680 210.000 ;
 END
END DOB37
PIN DIB36
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 993.920 208.880 995.040 210.000 ;
  LAYER metal4 ;
  RECT 993.920 208.880 995.040 210.000 ;
  LAYER metal3 ;
  RECT 993.920 208.880 995.040 210.000 ;
  LAYER metal2 ;
  RECT 993.920 208.880 995.040 210.000 ;
  LAYER metal1 ;
  RECT 993.920 208.880 995.040 210.000 ;
 END
END DIB36
PIN DOB36
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 980.280 208.880 981.400 210.000 ;
  LAYER metal4 ;
  RECT 980.280 208.880 981.400 210.000 ;
  LAYER metal3 ;
  RECT 980.280 208.880 981.400 210.000 ;
  LAYER metal2 ;
  RECT 980.280 208.880 981.400 210.000 ;
  LAYER metal1 ;
  RECT 980.280 208.880 981.400 210.000 ;
 END
END DOB36
PIN DIB35
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 967.260 208.880 968.380 210.000 ;
  LAYER metal4 ;
  RECT 967.260 208.880 968.380 210.000 ;
  LAYER metal3 ;
  RECT 967.260 208.880 968.380 210.000 ;
  LAYER metal2 ;
  RECT 967.260 208.880 968.380 210.000 ;
  LAYER metal1 ;
  RECT 967.260 208.880 968.380 210.000 ;
 END
END DIB35
PIN DOB35
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 953.620 208.880 954.740 210.000 ;
  LAYER metal4 ;
  RECT 953.620 208.880 954.740 210.000 ;
  LAYER metal3 ;
  RECT 953.620 208.880 954.740 210.000 ;
  LAYER metal2 ;
  RECT 953.620 208.880 954.740 210.000 ;
  LAYER metal1 ;
  RECT 953.620 208.880 954.740 210.000 ;
 END
END DOB35
PIN DIB34
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 939.980 208.880 941.100 210.000 ;
  LAYER metal4 ;
  RECT 939.980 208.880 941.100 210.000 ;
  LAYER metal3 ;
  RECT 939.980 208.880 941.100 210.000 ;
  LAYER metal2 ;
  RECT 939.980 208.880 941.100 210.000 ;
  LAYER metal1 ;
  RECT 939.980 208.880 941.100 210.000 ;
 END
END DIB34
PIN DOB34
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 926.960 208.880 928.080 210.000 ;
  LAYER metal4 ;
  RECT 926.960 208.880 928.080 210.000 ;
  LAYER metal3 ;
  RECT 926.960 208.880 928.080 210.000 ;
  LAYER metal2 ;
  RECT 926.960 208.880 928.080 210.000 ;
  LAYER metal1 ;
  RECT 926.960 208.880 928.080 210.000 ;
 END
END DOB34
PIN DIB33
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 913.320 208.880 914.440 210.000 ;
  LAYER metal4 ;
  RECT 913.320 208.880 914.440 210.000 ;
  LAYER metal3 ;
  RECT 913.320 208.880 914.440 210.000 ;
  LAYER metal2 ;
  RECT 913.320 208.880 914.440 210.000 ;
  LAYER metal1 ;
  RECT 913.320 208.880 914.440 210.000 ;
 END
END DIB33
PIN DOB33
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 899.680 208.880 900.800 210.000 ;
  LAYER metal4 ;
  RECT 899.680 208.880 900.800 210.000 ;
  LAYER metal3 ;
  RECT 899.680 208.880 900.800 210.000 ;
  LAYER metal2 ;
  RECT 899.680 208.880 900.800 210.000 ;
  LAYER metal1 ;
  RECT 899.680 208.880 900.800 210.000 ;
 END
END DOB33
PIN DIB32
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 886.040 208.880 887.160 210.000 ;
  LAYER metal4 ;
  RECT 886.040 208.880 887.160 210.000 ;
  LAYER metal3 ;
  RECT 886.040 208.880 887.160 210.000 ;
  LAYER metal2 ;
  RECT 886.040 208.880 887.160 210.000 ;
  LAYER metal1 ;
  RECT 886.040 208.880 887.160 210.000 ;
 END
END DIB32
PIN DOB32
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 873.020 208.880 874.140 210.000 ;
  LAYER metal4 ;
  RECT 873.020 208.880 874.140 210.000 ;
  LAYER metal3 ;
  RECT 873.020 208.880 874.140 210.000 ;
  LAYER metal2 ;
  RECT 873.020 208.880 874.140 210.000 ;
  LAYER metal1 ;
  RECT 873.020 208.880 874.140 210.000 ;
 END
END DOB32
PIN DIB31
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 859.380 208.880 860.500 210.000 ;
  LAYER metal4 ;
  RECT 859.380 208.880 860.500 210.000 ;
  LAYER metal3 ;
  RECT 859.380 208.880 860.500 210.000 ;
  LAYER metal2 ;
  RECT 859.380 208.880 860.500 210.000 ;
  LAYER metal1 ;
  RECT 859.380 208.880 860.500 210.000 ;
 END
END DIB31
PIN DOB31
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 845.740 208.880 846.860 210.000 ;
  LAYER metal4 ;
  RECT 845.740 208.880 846.860 210.000 ;
  LAYER metal3 ;
  RECT 845.740 208.880 846.860 210.000 ;
  LAYER metal2 ;
  RECT 845.740 208.880 846.860 210.000 ;
  LAYER metal1 ;
  RECT 845.740 208.880 846.860 210.000 ;
 END
END DOB31
PIN DIB30
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 832.720 208.880 833.840 210.000 ;
  LAYER metal4 ;
  RECT 832.720 208.880 833.840 210.000 ;
  LAYER metal3 ;
  RECT 832.720 208.880 833.840 210.000 ;
  LAYER metal2 ;
  RECT 832.720 208.880 833.840 210.000 ;
  LAYER metal1 ;
  RECT 832.720 208.880 833.840 210.000 ;
 END
END DIB30
PIN DOB30
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 819.080 208.880 820.200 210.000 ;
  LAYER metal4 ;
  RECT 819.080 208.880 820.200 210.000 ;
  LAYER metal3 ;
  RECT 819.080 208.880 820.200 210.000 ;
  LAYER metal2 ;
  RECT 819.080 208.880 820.200 210.000 ;
  LAYER metal1 ;
  RECT 819.080 208.880 820.200 210.000 ;
 END
END DOB30
PIN DIB29
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 805.440 208.880 806.560 210.000 ;
  LAYER metal4 ;
  RECT 805.440 208.880 806.560 210.000 ;
  LAYER metal3 ;
  RECT 805.440 208.880 806.560 210.000 ;
  LAYER metal2 ;
  RECT 805.440 208.880 806.560 210.000 ;
  LAYER metal1 ;
  RECT 805.440 208.880 806.560 210.000 ;
 END
END DIB29
PIN DOB29
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 792.420 208.880 793.540 210.000 ;
  LAYER metal4 ;
  RECT 792.420 208.880 793.540 210.000 ;
  LAYER metal3 ;
  RECT 792.420 208.880 793.540 210.000 ;
  LAYER metal2 ;
  RECT 792.420 208.880 793.540 210.000 ;
  LAYER metal1 ;
  RECT 792.420 208.880 793.540 210.000 ;
 END
END DOB29
PIN DIB28
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 778.780 208.880 779.900 210.000 ;
  LAYER metal4 ;
  RECT 778.780 208.880 779.900 210.000 ;
  LAYER metal3 ;
  RECT 778.780 208.880 779.900 210.000 ;
  LAYER metal2 ;
  RECT 778.780 208.880 779.900 210.000 ;
  LAYER metal1 ;
  RECT 778.780 208.880 779.900 210.000 ;
 END
END DIB28
PIN DOB28
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 765.140 208.880 766.260 210.000 ;
  LAYER metal4 ;
  RECT 765.140 208.880 766.260 210.000 ;
  LAYER metal3 ;
  RECT 765.140 208.880 766.260 210.000 ;
  LAYER metal2 ;
  RECT 765.140 208.880 766.260 210.000 ;
  LAYER metal1 ;
  RECT 765.140 208.880 766.260 210.000 ;
 END
END DOB28
PIN DIB27
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 752.120 208.880 753.240 210.000 ;
  LAYER metal4 ;
  RECT 752.120 208.880 753.240 210.000 ;
  LAYER metal3 ;
  RECT 752.120 208.880 753.240 210.000 ;
  LAYER metal2 ;
  RECT 752.120 208.880 753.240 210.000 ;
  LAYER metal1 ;
  RECT 752.120 208.880 753.240 210.000 ;
 END
END DIB27
PIN DOB27
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 738.480 208.880 739.600 210.000 ;
  LAYER metal4 ;
  RECT 738.480 208.880 739.600 210.000 ;
  LAYER metal3 ;
  RECT 738.480 208.880 739.600 210.000 ;
  LAYER metal2 ;
  RECT 738.480 208.880 739.600 210.000 ;
  LAYER metal1 ;
  RECT 738.480 208.880 739.600 210.000 ;
 END
END DOB27
PIN DIB26
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 724.840 208.880 725.960 210.000 ;
  LAYER metal4 ;
  RECT 724.840 208.880 725.960 210.000 ;
  LAYER metal3 ;
  RECT 724.840 208.880 725.960 210.000 ;
  LAYER metal2 ;
  RECT 724.840 208.880 725.960 210.000 ;
  LAYER metal1 ;
  RECT 724.840 208.880 725.960 210.000 ;
 END
END DIB26
PIN DOB26
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 711.820 208.880 712.940 210.000 ;
  LAYER metal4 ;
  RECT 711.820 208.880 712.940 210.000 ;
  LAYER metal3 ;
  RECT 711.820 208.880 712.940 210.000 ;
  LAYER metal2 ;
  RECT 711.820 208.880 712.940 210.000 ;
  LAYER metal1 ;
  RECT 711.820 208.880 712.940 210.000 ;
 END
END DOB26
PIN DIB25
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 698.180 208.880 699.300 210.000 ;
  LAYER metal4 ;
  RECT 698.180 208.880 699.300 210.000 ;
  LAYER metal3 ;
  RECT 698.180 208.880 699.300 210.000 ;
  LAYER metal2 ;
  RECT 698.180 208.880 699.300 210.000 ;
  LAYER metal1 ;
  RECT 698.180 208.880 699.300 210.000 ;
 END
END DIB25
PIN DOB25
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 684.540 208.880 685.660 210.000 ;
  LAYER metal4 ;
  RECT 684.540 208.880 685.660 210.000 ;
  LAYER metal3 ;
  RECT 684.540 208.880 685.660 210.000 ;
  LAYER metal2 ;
  RECT 684.540 208.880 685.660 210.000 ;
  LAYER metal1 ;
  RECT 684.540 208.880 685.660 210.000 ;
 END
END DOB25
PIN DIB24
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 671.520 208.880 672.640 210.000 ;
  LAYER metal4 ;
  RECT 671.520 208.880 672.640 210.000 ;
  LAYER metal3 ;
  RECT 671.520 208.880 672.640 210.000 ;
  LAYER metal2 ;
  RECT 671.520 208.880 672.640 210.000 ;
  LAYER metal1 ;
  RECT 671.520 208.880 672.640 210.000 ;
 END
END DIB24
PIN DOB24
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 657.880 208.880 659.000 210.000 ;
  LAYER metal4 ;
  RECT 657.880 208.880 659.000 210.000 ;
  LAYER metal3 ;
  RECT 657.880 208.880 659.000 210.000 ;
  LAYER metal2 ;
  RECT 657.880 208.880 659.000 210.000 ;
  LAYER metal1 ;
  RECT 657.880 208.880 659.000 210.000 ;
 END
END DOB24
PIN DIB23
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 644.240 208.880 645.360 210.000 ;
  LAYER metal4 ;
  RECT 644.240 208.880 645.360 210.000 ;
  LAYER metal3 ;
  RECT 644.240 208.880 645.360 210.000 ;
  LAYER metal2 ;
  RECT 644.240 208.880 645.360 210.000 ;
  LAYER metal1 ;
  RECT 644.240 208.880 645.360 210.000 ;
 END
END DIB23
PIN DOB23
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 631.220 208.880 632.340 210.000 ;
  LAYER metal4 ;
  RECT 631.220 208.880 632.340 210.000 ;
  LAYER metal3 ;
  RECT 631.220 208.880 632.340 210.000 ;
  LAYER metal2 ;
  RECT 631.220 208.880 632.340 210.000 ;
  LAYER metal1 ;
  RECT 631.220 208.880 632.340 210.000 ;
 END
END DOB23
PIN DIB22
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 617.580 208.880 618.700 210.000 ;
  LAYER metal4 ;
  RECT 617.580 208.880 618.700 210.000 ;
  LAYER metal3 ;
  RECT 617.580 208.880 618.700 210.000 ;
  LAYER metal2 ;
  RECT 617.580 208.880 618.700 210.000 ;
  LAYER metal1 ;
  RECT 617.580 208.880 618.700 210.000 ;
 END
END DIB22
PIN DOB22
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 603.940 208.880 605.060 210.000 ;
  LAYER metal4 ;
  RECT 603.940 208.880 605.060 210.000 ;
  LAYER metal3 ;
  RECT 603.940 208.880 605.060 210.000 ;
  LAYER metal2 ;
  RECT 603.940 208.880 605.060 210.000 ;
  LAYER metal1 ;
  RECT 603.940 208.880 605.060 210.000 ;
 END
END DOB22
PIN DIB21
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 590.920 208.880 592.040 210.000 ;
  LAYER metal4 ;
  RECT 590.920 208.880 592.040 210.000 ;
  LAYER metal3 ;
  RECT 590.920 208.880 592.040 210.000 ;
  LAYER metal2 ;
  RECT 590.920 208.880 592.040 210.000 ;
  LAYER metal1 ;
  RECT 590.920 208.880 592.040 210.000 ;
 END
END DIB21
PIN DOB21
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 577.280 208.880 578.400 210.000 ;
  LAYER metal4 ;
  RECT 577.280 208.880 578.400 210.000 ;
  LAYER metal3 ;
  RECT 577.280 208.880 578.400 210.000 ;
  LAYER metal2 ;
  RECT 577.280 208.880 578.400 210.000 ;
  LAYER metal1 ;
  RECT 577.280 208.880 578.400 210.000 ;
 END
END DOB21
PIN DIB20
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 563.640 208.880 564.760 210.000 ;
  LAYER metal4 ;
  RECT 563.640 208.880 564.760 210.000 ;
  LAYER metal3 ;
  RECT 563.640 208.880 564.760 210.000 ;
  LAYER metal2 ;
  RECT 563.640 208.880 564.760 210.000 ;
  LAYER metal1 ;
  RECT 563.640 208.880 564.760 210.000 ;
 END
END DIB20
PIN DOB20
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 550.620 208.880 551.740 210.000 ;
  LAYER metal4 ;
  RECT 550.620 208.880 551.740 210.000 ;
  LAYER metal3 ;
  RECT 550.620 208.880 551.740 210.000 ;
  LAYER metal2 ;
  RECT 550.620 208.880 551.740 210.000 ;
  LAYER metal1 ;
  RECT 550.620 208.880 551.740 210.000 ;
 END
END DOB20
PIN DIB19
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 536.980 208.880 538.100 210.000 ;
  LAYER metal4 ;
  RECT 536.980 208.880 538.100 210.000 ;
  LAYER metal3 ;
  RECT 536.980 208.880 538.100 210.000 ;
  LAYER metal2 ;
  RECT 536.980 208.880 538.100 210.000 ;
  LAYER metal1 ;
  RECT 536.980 208.880 538.100 210.000 ;
 END
END DIB19
PIN DOB19
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 523.340 208.880 524.460 210.000 ;
  LAYER metal4 ;
  RECT 523.340 208.880 524.460 210.000 ;
  LAYER metal3 ;
  RECT 523.340 208.880 524.460 210.000 ;
  LAYER metal2 ;
  RECT 523.340 208.880 524.460 210.000 ;
  LAYER metal1 ;
  RECT 523.340 208.880 524.460 210.000 ;
 END
END DOB19
PIN DIB18
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 510.320 208.880 511.440 210.000 ;
  LAYER metal4 ;
  RECT 510.320 208.880 511.440 210.000 ;
  LAYER metal3 ;
  RECT 510.320 208.880 511.440 210.000 ;
  LAYER metal2 ;
  RECT 510.320 208.880 511.440 210.000 ;
  LAYER metal1 ;
  RECT 510.320 208.880 511.440 210.000 ;
 END
END DIB18
PIN DOB18
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 496.680 208.880 497.800 210.000 ;
  LAYER metal4 ;
  RECT 496.680 208.880 497.800 210.000 ;
  LAYER metal3 ;
  RECT 496.680 208.880 497.800 210.000 ;
  LAYER metal2 ;
  RECT 496.680 208.880 497.800 210.000 ;
  LAYER metal1 ;
  RECT 496.680 208.880 497.800 210.000 ;
 END
END DOB18
PIN DIB17
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 483.040 208.880 484.160 210.000 ;
  LAYER metal4 ;
  RECT 483.040 208.880 484.160 210.000 ;
  LAYER metal3 ;
  RECT 483.040 208.880 484.160 210.000 ;
  LAYER metal2 ;
  RECT 483.040 208.880 484.160 210.000 ;
  LAYER metal1 ;
  RECT 483.040 208.880 484.160 210.000 ;
 END
END DIB17
PIN DOB17
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 469.400 208.880 470.520 210.000 ;
  LAYER metal4 ;
  RECT 469.400 208.880 470.520 210.000 ;
  LAYER metal3 ;
  RECT 469.400 208.880 470.520 210.000 ;
  LAYER metal2 ;
  RECT 469.400 208.880 470.520 210.000 ;
  LAYER metal1 ;
  RECT 469.400 208.880 470.520 210.000 ;
 END
END DOB17
PIN DIB16
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 456.380 208.880 457.500 210.000 ;
  LAYER metal4 ;
  RECT 456.380 208.880 457.500 210.000 ;
  LAYER metal3 ;
  RECT 456.380 208.880 457.500 210.000 ;
  LAYER metal2 ;
  RECT 456.380 208.880 457.500 210.000 ;
  LAYER metal1 ;
  RECT 456.380 208.880 457.500 210.000 ;
 END
END DIB16
PIN DOB16
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 442.740 208.880 443.860 210.000 ;
  LAYER metal4 ;
  RECT 442.740 208.880 443.860 210.000 ;
  LAYER metal3 ;
  RECT 442.740 208.880 443.860 210.000 ;
  LAYER metal2 ;
  RECT 442.740 208.880 443.860 210.000 ;
  LAYER metal1 ;
  RECT 442.740 208.880 443.860 210.000 ;
 END
END DOB16
PIN DIB15
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 429.100 208.880 430.220 210.000 ;
  LAYER metal4 ;
  RECT 429.100 208.880 430.220 210.000 ;
  LAYER metal3 ;
  RECT 429.100 208.880 430.220 210.000 ;
  LAYER metal2 ;
  RECT 429.100 208.880 430.220 210.000 ;
  LAYER metal1 ;
  RECT 429.100 208.880 430.220 210.000 ;
 END
END DIB15
PIN DOB15
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 416.080 208.880 417.200 210.000 ;
  LAYER metal4 ;
  RECT 416.080 208.880 417.200 210.000 ;
  LAYER metal3 ;
  RECT 416.080 208.880 417.200 210.000 ;
  LAYER metal2 ;
  RECT 416.080 208.880 417.200 210.000 ;
  LAYER metal1 ;
  RECT 416.080 208.880 417.200 210.000 ;
 END
END DOB15
PIN DIB14
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 402.440 208.880 403.560 210.000 ;
  LAYER metal4 ;
  RECT 402.440 208.880 403.560 210.000 ;
  LAYER metal3 ;
  RECT 402.440 208.880 403.560 210.000 ;
  LAYER metal2 ;
  RECT 402.440 208.880 403.560 210.000 ;
  LAYER metal1 ;
  RECT 402.440 208.880 403.560 210.000 ;
 END
END DIB14
PIN DOB14
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 388.800 208.880 389.920 210.000 ;
  LAYER metal4 ;
  RECT 388.800 208.880 389.920 210.000 ;
  LAYER metal3 ;
  RECT 388.800 208.880 389.920 210.000 ;
  LAYER metal2 ;
  RECT 388.800 208.880 389.920 210.000 ;
  LAYER metal1 ;
  RECT 388.800 208.880 389.920 210.000 ;
 END
END DOB14
PIN DIB13
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 375.780 208.880 376.900 210.000 ;
  LAYER metal4 ;
  RECT 375.780 208.880 376.900 210.000 ;
  LAYER metal3 ;
  RECT 375.780 208.880 376.900 210.000 ;
  LAYER metal2 ;
  RECT 375.780 208.880 376.900 210.000 ;
  LAYER metal1 ;
  RECT 375.780 208.880 376.900 210.000 ;
 END
END DIB13
PIN DOB13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 362.140 208.880 363.260 210.000 ;
  LAYER metal4 ;
  RECT 362.140 208.880 363.260 210.000 ;
  LAYER metal3 ;
  RECT 362.140 208.880 363.260 210.000 ;
  LAYER metal2 ;
  RECT 362.140 208.880 363.260 210.000 ;
  LAYER metal1 ;
  RECT 362.140 208.880 363.260 210.000 ;
 END
END DOB13
PIN DIB12
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 348.500 208.880 349.620 210.000 ;
  LAYER metal4 ;
  RECT 348.500 208.880 349.620 210.000 ;
  LAYER metal3 ;
  RECT 348.500 208.880 349.620 210.000 ;
  LAYER metal2 ;
  RECT 348.500 208.880 349.620 210.000 ;
  LAYER metal1 ;
  RECT 348.500 208.880 349.620 210.000 ;
 END
END DIB12
PIN DOB12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 335.480 208.880 336.600 210.000 ;
  LAYER metal4 ;
  RECT 335.480 208.880 336.600 210.000 ;
  LAYER metal3 ;
  RECT 335.480 208.880 336.600 210.000 ;
  LAYER metal2 ;
  RECT 335.480 208.880 336.600 210.000 ;
  LAYER metal1 ;
  RECT 335.480 208.880 336.600 210.000 ;
 END
END DOB12
PIN DIB11
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 321.840 208.880 322.960 210.000 ;
  LAYER metal4 ;
  RECT 321.840 208.880 322.960 210.000 ;
  LAYER metal3 ;
  RECT 321.840 208.880 322.960 210.000 ;
  LAYER metal2 ;
  RECT 321.840 208.880 322.960 210.000 ;
  LAYER metal1 ;
  RECT 321.840 208.880 322.960 210.000 ;
 END
END DIB11
PIN DOB11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 308.200 208.880 309.320 210.000 ;
  LAYER metal4 ;
  RECT 308.200 208.880 309.320 210.000 ;
  LAYER metal3 ;
  RECT 308.200 208.880 309.320 210.000 ;
  LAYER metal2 ;
  RECT 308.200 208.880 309.320 210.000 ;
  LAYER metal1 ;
  RECT 308.200 208.880 309.320 210.000 ;
 END
END DOB11
PIN DIB10
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 295.180 208.880 296.300 210.000 ;
  LAYER metal4 ;
  RECT 295.180 208.880 296.300 210.000 ;
  LAYER metal3 ;
  RECT 295.180 208.880 296.300 210.000 ;
  LAYER metal2 ;
  RECT 295.180 208.880 296.300 210.000 ;
  LAYER metal1 ;
  RECT 295.180 208.880 296.300 210.000 ;
 END
END DIB10
PIN DOB10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 281.540 208.880 282.660 210.000 ;
  LAYER metal4 ;
  RECT 281.540 208.880 282.660 210.000 ;
  LAYER metal3 ;
  RECT 281.540 208.880 282.660 210.000 ;
  LAYER metal2 ;
  RECT 281.540 208.880 282.660 210.000 ;
  LAYER metal1 ;
  RECT 281.540 208.880 282.660 210.000 ;
 END
END DOB10
PIN DIB9
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 267.900 208.880 269.020 210.000 ;
  LAYER metal4 ;
  RECT 267.900 208.880 269.020 210.000 ;
  LAYER metal3 ;
  RECT 267.900 208.880 269.020 210.000 ;
  LAYER metal2 ;
  RECT 267.900 208.880 269.020 210.000 ;
  LAYER metal1 ;
  RECT 267.900 208.880 269.020 210.000 ;
 END
END DIB9
PIN DOB9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 254.880 208.880 256.000 210.000 ;
  LAYER metal4 ;
  RECT 254.880 208.880 256.000 210.000 ;
  LAYER metal3 ;
  RECT 254.880 208.880 256.000 210.000 ;
  LAYER metal2 ;
  RECT 254.880 208.880 256.000 210.000 ;
  LAYER metal1 ;
  RECT 254.880 208.880 256.000 210.000 ;
 END
END DOB9
PIN DIB8
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 241.240 208.880 242.360 210.000 ;
  LAYER metal4 ;
  RECT 241.240 208.880 242.360 210.000 ;
  LAYER metal3 ;
  RECT 241.240 208.880 242.360 210.000 ;
  LAYER metal2 ;
  RECT 241.240 208.880 242.360 210.000 ;
  LAYER metal1 ;
  RECT 241.240 208.880 242.360 210.000 ;
 END
END DIB8
PIN DOB8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 227.600 208.880 228.720 210.000 ;
  LAYER metal4 ;
  RECT 227.600 208.880 228.720 210.000 ;
  LAYER metal3 ;
  RECT 227.600 208.880 228.720 210.000 ;
  LAYER metal2 ;
  RECT 227.600 208.880 228.720 210.000 ;
  LAYER metal1 ;
  RECT 227.600 208.880 228.720 210.000 ;
 END
END DOB8
PIN DIB7
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 214.580 208.880 215.700 210.000 ;
  LAYER metal4 ;
  RECT 214.580 208.880 215.700 210.000 ;
  LAYER metal3 ;
  RECT 214.580 208.880 215.700 210.000 ;
  LAYER metal2 ;
  RECT 214.580 208.880 215.700 210.000 ;
  LAYER metal1 ;
  RECT 214.580 208.880 215.700 210.000 ;
 END
END DIB7
PIN DOB7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 200.940 208.880 202.060 210.000 ;
  LAYER metal4 ;
  RECT 200.940 208.880 202.060 210.000 ;
  LAYER metal3 ;
  RECT 200.940 208.880 202.060 210.000 ;
  LAYER metal2 ;
  RECT 200.940 208.880 202.060 210.000 ;
  LAYER metal1 ;
  RECT 200.940 208.880 202.060 210.000 ;
 END
END DOB7
PIN DIB6
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 187.300 208.880 188.420 210.000 ;
  LAYER metal4 ;
  RECT 187.300 208.880 188.420 210.000 ;
  LAYER metal3 ;
  RECT 187.300 208.880 188.420 210.000 ;
  LAYER metal2 ;
  RECT 187.300 208.880 188.420 210.000 ;
  LAYER metal1 ;
  RECT 187.300 208.880 188.420 210.000 ;
 END
END DIB6
PIN DOB6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 174.280 208.880 175.400 210.000 ;
  LAYER metal4 ;
  RECT 174.280 208.880 175.400 210.000 ;
  LAYER metal3 ;
  RECT 174.280 208.880 175.400 210.000 ;
  LAYER metal2 ;
  RECT 174.280 208.880 175.400 210.000 ;
  LAYER metal1 ;
  RECT 174.280 208.880 175.400 210.000 ;
 END
END DOB6
PIN DIB5
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 160.640 208.880 161.760 210.000 ;
  LAYER metal4 ;
  RECT 160.640 208.880 161.760 210.000 ;
  LAYER metal3 ;
  RECT 160.640 208.880 161.760 210.000 ;
  LAYER metal2 ;
  RECT 160.640 208.880 161.760 210.000 ;
  LAYER metal1 ;
  RECT 160.640 208.880 161.760 210.000 ;
 END
END DIB5
PIN DOB5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 147.000 208.880 148.120 210.000 ;
  LAYER metal4 ;
  RECT 147.000 208.880 148.120 210.000 ;
  LAYER metal3 ;
  RECT 147.000 208.880 148.120 210.000 ;
  LAYER metal2 ;
  RECT 147.000 208.880 148.120 210.000 ;
  LAYER metal1 ;
  RECT 147.000 208.880 148.120 210.000 ;
 END
END DOB5
PIN DIB4
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 133.980 208.880 135.100 210.000 ;
  LAYER metal4 ;
  RECT 133.980 208.880 135.100 210.000 ;
  LAYER metal3 ;
  RECT 133.980 208.880 135.100 210.000 ;
  LAYER metal2 ;
  RECT 133.980 208.880 135.100 210.000 ;
  LAYER metal1 ;
  RECT 133.980 208.880 135.100 210.000 ;
 END
END DIB4
PIN DOB4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 120.340 208.880 121.460 210.000 ;
  LAYER metal4 ;
  RECT 120.340 208.880 121.460 210.000 ;
  LAYER metal3 ;
  RECT 120.340 208.880 121.460 210.000 ;
  LAYER metal2 ;
  RECT 120.340 208.880 121.460 210.000 ;
  LAYER metal1 ;
  RECT 120.340 208.880 121.460 210.000 ;
 END
END DOB4
PIN DIB3
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 106.700 208.880 107.820 210.000 ;
  LAYER metal4 ;
  RECT 106.700 208.880 107.820 210.000 ;
  LAYER metal3 ;
  RECT 106.700 208.880 107.820 210.000 ;
  LAYER metal2 ;
  RECT 106.700 208.880 107.820 210.000 ;
  LAYER metal1 ;
  RECT 106.700 208.880 107.820 210.000 ;
 END
END DIB3
PIN DOB3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 93.680 208.880 94.800 210.000 ;
  LAYER metal4 ;
  RECT 93.680 208.880 94.800 210.000 ;
  LAYER metal3 ;
  RECT 93.680 208.880 94.800 210.000 ;
  LAYER metal2 ;
  RECT 93.680 208.880 94.800 210.000 ;
  LAYER metal1 ;
  RECT 93.680 208.880 94.800 210.000 ;
 END
END DOB3
PIN DIB2
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 80.040 208.880 81.160 210.000 ;
  LAYER metal4 ;
  RECT 80.040 208.880 81.160 210.000 ;
  LAYER metal3 ;
  RECT 80.040 208.880 81.160 210.000 ;
  LAYER metal2 ;
  RECT 80.040 208.880 81.160 210.000 ;
  LAYER metal1 ;
  RECT 80.040 208.880 81.160 210.000 ;
 END
END DIB2
PIN DOB2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 66.400 208.880 67.520 210.000 ;
  LAYER metal4 ;
  RECT 66.400 208.880 67.520 210.000 ;
  LAYER metal3 ;
  RECT 66.400 208.880 67.520 210.000 ;
  LAYER metal2 ;
  RECT 66.400 208.880 67.520 210.000 ;
  LAYER metal1 ;
  RECT 66.400 208.880 67.520 210.000 ;
 END
END DOB2
PIN DIB1
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 52.760 208.880 53.880 210.000 ;
  LAYER metal4 ;
  RECT 52.760 208.880 53.880 210.000 ;
  LAYER metal3 ;
  RECT 52.760 208.880 53.880 210.000 ;
  LAYER metal2 ;
  RECT 52.760 208.880 53.880 210.000 ;
  LAYER metal1 ;
  RECT 52.760 208.880 53.880 210.000 ;
 END
END DIB1
PIN DOB1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 39.740 208.880 40.860 210.000 ;
  LAYER metal4 ;
  RECT 39.740 208.880 40.860 210.000 ;
  LAYER metal3 ;
  RECT 39.740 208.880 40.860 210.000 ;
  LAYER metal2 ;
  RECT 39.740 208.880 40.860 210.000 ;
  LAYER metal1 ;
  RECT 39.740 208.880 40.860 210.000 ;
 END
END DOB1
PIN DIB0
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 26.100 208.880 27.220 210.000 ;
  LAYER metal4 ;
  RECT 26.100 208.880 27.220 210.000 ;
  LAYER metal3 ;
  RECT 26.100 208.880 27.220 210.000 ;
  LAYER metal2 ;
  RECT 26.100 208.880 27.220 210.000 ;
  LAYER metal1 ;
  RECT 26.100 208.880 27.220 210.000 ;
 END
END DIB0
PIN DOB0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 12.460 208.880 13.580 210.000 ;
  LAYER metal4 ;
  RECT 12.460 208.880 13.580 210.000 ;
  LAYER metal3 ;
  RECT 12.460 208.880 13.580 210.000 ;
  LAYER metal2 ;
  RECT 12.460 208.880 13.580 210.000 ;
  LAYER metal1 ;
  RECT 12.460 208.880 13.580 210.000 ;
 END
END DOB0
PIN DIA127
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3548.940 0.000 3550.060 1.120 ;
  LAYER metal4 ;
  RECT 3548.940 0.000 3550.060 1.120 ;
  LAYER metal3 ;
  RECT 3548.940 0.000 3550.060 1.120 ;
  LAYER metal2 ;
  RECT 3548.940 0.000 3550.060 1.120 ;
  LAYER metal1 ;
  RECT 3548.940 0.000 3550.060 1.120 ;
 END
END DIA127
PIN DOA127
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3535.300 0.000 3536.420 1.120 ;
  LAYER metal4 ;
  RECT 3535.300 0.000 3536.420 1.120 ;
  LAYER metal3 ;
  RECT 3535.300 0.000 3536.420 1.120 ;
  LAYER metal2 ;
  RECT 3535.300 0.000 3536.420 1.120 ;
  LAYER metal1 ;
  RECT 3535.300 0.000 3536.420 1.120 ;
 END
END DOA127
PIN DIA126
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3522.280 0.000 3523.400 1.120 ;
  LAYER metal4 ;
  RECT 3522.280 0.000 3523.400 1.120 ;
  LAYER metal3 ;
  RECT 3522.280 0.000 3523.400 1.120 ;
  LAYER metal2 ;
  RECT 3522.280 0.000 3523.400 1.120 ;
  LAYER metal1 ;
  RECT 3522.280 0.000 3523.400 1.120 ;
 END
END DIA126
PIN DOA126
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3508.640 0.000 3509.760 1.120 ;
  LAYER metal4 ;
  RECT 3508.640 0.000 3509.760 1.120 ;
  LAYER metal3 ;
  RECT 3508.640 0.000 3509.760 1.120 ;
  LAYER metal2 ;
  RECT 3508.640 0.000 3509.760 1.120 ;
  LAYER metal1 ;
  RECT 3508.640 0.000 3509.760 1.120 ;
 END
END DOA126
PIN DIA125
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3495.000 0.000 3496.120 1.120 ;
  LAYER metal4 ;
  RECT 3495.000 0.000 3496.120 1.120 ;
  LAYER metal3 ;
  RECT 3495.000 0.000 3496.120 1.120 ;
  LAYER metal2 ;
  RECT 3495.000 0.000 3496.120 1.120 ;
  LAYER metal1 ;
  RECT 3495.000 0.000 3496.120 1.120 ;
 END
END DIA125
PIN DOA125
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3481.980 0.000 3483.100 1.120 ;
  LAYER metal4 ;
  RECT 3481.980 0.000 3483.100 1.120 ;
  LAYER metal3 ;
  RECT 3481.980 0.000 3483.100 1.120 ;
  LAYER metal2 ;
  RECT 3481.980 0.000 3483.100 1.120 ;
  LAYER metal1 ;
  RECT 3481.980 0.000 3483.100 1.120 ;
 END
END DOA125
PIN DIA124
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3468.340 0.000 3469.460 1.120 ;
  LAYER metal4 ;
  RECT 3468.340 0.000 3469.460 1.120 ;
  LAYER metal3 ;
  RECT 3468.340 0.000 3469.460 1.120 ;
  LAYER metal2 ;
  RECT 3468.340 0.000 3469.460 1.120 ;
  LAYER metal1 ;
  RECT 3468.340 0.000 3469.460 1.120 ;
 END
END DIA124
PIN DOA124
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3454.700 0.000 3455.820 1.120 ;
  LAYER metal4 ;
  RECT 3454.700 0.000 3455.820 1.120 ;
  LAYER metal3 ;
  RECT 3454.700 0.000 3455.820 1.120 ;
  LAYER metal2 ;
  RECT 3454.700 0.000 3455.820 1.120 ;
  LAYER metal1 ;
  RECT 3454.700 0.000 3455.820 1.120 ;
 END
END DOA124
PIN DIA123
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3441.060 0.000 3442.180 1.120 ;
  LAYER metal4 ;
  RECT 3441.060 0.000 3442.180 1.120 ;
  LAYER metal3 ;
  RECT 3441.060 0.000 3442.180 1.120 ;
  LAYER metal2 ;
  RECT 3441.060 0.000 3442.180 1.120 ;
  LAYER metal1 ;
  RECT 3441.060 0.000 3442.180 1.120 ;
 END
END DIA123
PIN DOA123
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3428.040 0.000 3429.160 1.120 ;
  LAYER metal4 ;
  RECT 3428.040 0.000 3429.160 1.120 ;
  LAYER metal3 ;
  RECT 3428.040 0.000 3429.160 1.120 ;
  LAYER metal2 ;
  RECT 3428.040 0.000 3429.160 1.120 ;
  LAYER metal1 ;
  RECT 3428.040 0.000 3429.160 1.120 ;
 END
END DOA123
PIN DIA122
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3414.400 0.000 3415.520 1.120 ;
  LAYER metal4 ;
  RECT 3414.400 0.000 3415.520 1.120 ;
  LAYER metal3 ;
  RECT 3414.400 0.000 3415.520 1.120 ;
  LAYER metal2 ;
  RECT 3414.400 0.000 3415.520 1.120 ;
  LAYER metal1 ;
  RECT 3414.400 0.000 3415.520 1.120 ;
 END
END DIA122
PIN DOA122
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3400.760 0.000 3401.880 1.120 ;
  LAYER metal4 ;
  RECT 3400.760 0.000 3401.880 1.120 ;
  LAYER metal3 ;
  RECT 3400.760 0.000 3401.880 1.120 ;
  LAYER metal2 ;
  RECT 3400.760 0.000 3401.880 1.120 ;
  LAYER metal1 ;
  RECT 3400.760 0.000 3401.880 1.120 ;
 END
END DOA122
PIN DIA121
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3387.740 0.000 3388.860 1.120 ;
  LAYER metal4 ;
  RECT 3387.740 0.000 3388.860 1.120 ;
  LAYER metal3 ;
  RECT 3387.740 0.000 3388.860 1.120 ;
  LAYER metal2 ;
  RECT 3387.740 0.000 3388.860 1.120 ;
  LAYER metal1 ;
  RECT 3387.740 0.000 3388.860 1.120 ;
 END
END DIA121
PIN DOA121
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3374.100 0.000 3375.220 1.120 ;
  LAYER metal4 ;
  RECT 3374.100 0.000 3375.220 1.120 ;
  LAYER metal3 ;
  RECT 3374.100 0.000 3375.220 1.120 ;
  LAYER metal2 ;
  RECT 3374.100 0.000 3375.220 1.120 ;
  LAYER metal1 ;
  RECT 3374.100 0.000 3375.220 1.120 ;
 END
END DOA121
PIN DIA120
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3360.460 0.000 3361.580 1.120 ;
  LAYER metal4 ;
  RECT 3360.460 0.000 3361.580 1.120 ;
  LAYER metal3 ;
  RECT 3360.460 0.000 3361.580 1.120 ;
  LAYER metal2 ;
  RECT 3360.460 0.000 3361.580 1.120 ;
  LAYER metal1 ;
  RECT 3360.460 0.000 3361.580 1.120 ;
 END
END DIA120
PIN DOA120
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3347.440 0.000 3348.560 1.120 ;
  LAYER metal4 ;
  RECT 3347.440 0.000 3348.560 1.120 ;
  LAYER metal3 ;
  RECT 3347.440 0.000 3348.560 1.120 ;
  LAYER metal2 ;
  RECT 3347.440 0.000 3348.560 1.120 ;
  LAYER metal1 ;
  RECT 3347.440 0.000 3348.560 1.120 ;
 END
END DOA120
PIN DIA119
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3333.800 0.000 3334.920 1.120 ;
  LAYER metal4 ;
  RECT 3333.800 0.000 3334.920 1.120 ;
  LAYER metal3 ;
  RECT 3333.800 0.000 3334.920 1.120 ;
  LAYER metal2 ;
  RECT 3333.800 0.000 3334.920 1.120 ;
  LAYER metal1 ;
  RECT 3333.800 0.000 3334.920 1.120 ;
 END
END DIA119
PIN DOA119
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3320.160 0.000 3321.280 1.120 ;
  LAYER metal4 ;
  RECT 3320.160 0.000 3321.280 1.120 ;
  LAYER metal3 ;
  RECT 3320.160 0.000 3321.280 1.120 ;
  LAYER metal2 ;
  RECT 3320.160 0.000 3321.280 1.120 ;
  LAYER metal1 ;
  RECT 3320.160 0.000 3321.280 1.120 ;
 END
END DOA119
PIN DIA118
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3307.140 0.000 3308.260 1.120 ;
  LAYER metal4 ;
  RECT 3307.140 0.000 3308.260 1.120 ;
  LAYER metal3 ;
  RECT 3307.140 0.000 3308.260 1.120 ;
  LAYER metal2 ;
  RECT 3307.140 0.000 3308.260 1.120 ;
  LAYER metal1 ;
  RECT 3307.140 0.000 3308.260 1.120 ;
 END
END DIA118
PIN DOA118
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3293.500 0.000 3294.620 1.120 ;
  LAYER metal4 ;
  RECT 3293.500 0.000 3294.620 1.120 ;
  LAYER metal3 ;
  RECT 3293.500 0.000 3294.620 1.120 ;
  LAYER metal2 ;
  RECT 3293.500 0.000 3294.620 1.120 ;
  LAYER metal1 ;
  RECT 3293.500 0.000 3294.620 1.120 ;
 END
END DOA118
PIN DIA117
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3279.860 0.000 3280.980 1.120 ;
  LAYER metal4 ;
  RECT 3279.860 0.000 3280.980 1.120 ;
  LAYER metal3 ;
  RECT 3279.860 0.000 3280.980 1.120 ;
  LAYER metal2 ;
  RECT 3279.860 0.000 3280.980 1.120 ;
  LAYER metal1 ;
  RECT 3279.860 0.000 3280.980 1.120 ;
 END
END DIA117
PIN DOA117
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3266.840 0.000 3267.960 1.120 ;
  LAYER metal4 ;
  RECT 3266.840 0.000 3267.960 1.120 ;
  LAYER metal3 ;
  RECT 3266.840 0.000 3267.960 1.120 ;
  LAYER metal2 ;
  RECT 3266.840 0.000 3267.960 1.120 ;
  LAYER metal1 ;
  RECT 3266.840 0.000 3267.960 1.120 ;
 END
END DOA117
PIN DIA116
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3253.200 0.000 3254.320 1.120 ;
  LAYER metal4 ;
  RECT 3253.200 0.000 3254.320 1.120 ;
  LAYER metal3 ;
  RECT 3253.200 0.000 3254.320 1.120 ;
  LAYER metal2 ;
  RECT 3253.200 0.000 3254.320 1.120 ;
  LAYER metal1 ;
  RECT 3253.200 0.000 3254.320 1.120 ;
 END
END DIA116
PIN DOA116
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3239.560 0.000 3240.680 1.120 ;
  LAYER metal4 ;
  RECT 3239.560 0.000 3240.680 1.120 ;
  LAYER metal3 ;
  RECT 3239.560 0.000 3240.680 1.120 ;
  LAYER metal2 ;
  RECT 3239.560 0.000 3240.680 1.120 ;
  LAYER metal1 ;
  RECT 3239.560 0.000 3240.680 1.120 ;
 END
END DOA116
PIN DIA115
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3226.540 0.000 3227.660 1.120 ;
  LAYER metal4 ;
  RECT 3226.540 0.000 3227.660 1.120 ;
  LAYER metal3 ;
  RECT 3226.540 0.000 3227.660 1.120 ;
  LAYER metal2 ;
  RECT 3226.540 0.000 3227.660 1.120 ;
  LAYER metal1 ;
  RECT 3226.540 0.000 3227.660 1.120 ;
 END
END DIA115
PIN DOA115
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3212.900 0.000 3214.020 1.120 ;
  LAYER metal4 ;
  RECT 3212.900 0.000 3214.020 1.120 ;
  LAYER metal3 ;
  RECT 3212.900 0.000 3214.020 1.120 ;
  LAYER metal2 ;
  RECT 3212.900 0.000 3214.020 1.120 ;
  LAYER metal1 ;
  RECT 3212.900 0.000 3214.020 1.120 ;
 END
END DOA115
PIN DIA114
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3199.260 0.000 3200.380 1.120 ;
  LAYER metal4 ;
  RECT 3199.260 0.000 3200.380 1.120 ;
  LAYER metal3 ;
  RECT 3199.260 0.000 3200.380 1.120 ;
  LAYER metal2 ;
  RECT 3199.260 0.000 3200.380 1.120 ;
  LAYER metal1 ;
  RECT 3199.260 0.000 3200.380 1.120 ;
 END
END DIA114
PIN DOA114
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3186.240 0.000 3187.360 1.120 ;
  LAYER metal4 ;
  RECT 3186.240 0.000 3187.360 1.120 ;
  LAYER metal3 ;
  RECT 3186.240 0.000 3187.360 1.120 ;
  LAYER metal2 ;
  RECT 3186.240 0.000 3187.360 1.120 ;
  LAYER metal1 ;
  RECT 3186.240 0.000 3187.360 1.120 ;
 END
END DOA114
PIN DIA113
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3172.600 0.000 3173.720 1.120 ;
  LAYER metal4 ;
  RECT 3172.600 0.000 3173.720 1.120 ;
  LAYER metal3 ;
  RECT 3172.600 0.000 3173.720 1.120 ;
  LAYER metal2 ;
  RECT 3172.600 0.000 3173.720 1.120 ;
  LAYER metal1 ;
  RECT 3172.600 0.000 3173.720 1.120 ;
 END
END DIA113
PIN DOA113
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3158.960 0.000 3160.080 1.120 ;
  LAYER metal4 ;
  RECT 3158.960 0.000 3160.080 1.120 ;
  LAYER metal3 ;
  RECT 3158.960 0.000 3160.080 1.120 ;
  LAYER metal2 ;
  RECT 3158.960 0.000 3160.080 1.120 ;
  LAYER metal1 ;
  RECT 3158.960 0.000 3160.080 1.120 ;
 END
END DOA113
PIN DIA112
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3145.940 0.000 3147.060 1.120 ;
  LAYER metal4 ;
  RECT 3145.940 0.000 3147.060 1.120 ;
  LAYER metal3 ;
  RECT 3145.940 0.000 3147.060 1.120 ;
  LAYER metal2 ;
  RECT 3145.940 0.000 3147.060 1.120 ;
  LAYER metal1 ;
  RECT 3145.940 0.000 3147.060 1.120 ;
 END
END DIA112
PIN DOA112
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3132.300 0.000 3133.420 1.120 ;
  LAYER metal4 ;
  RECT 3132.300 0.000 3133.420 1.120 ;
  LAYER metal3 ;
  RECT 3132.300 0.000 3133.420 1.120 ;
  LAYER metal2 ;
  RECT 3132.300 0.000 3133.420 1.120 ;
  LAYER metal1 ;
  RECT 3132.300 0.000 3133.420 1.120 ;
 END
END DOA112
PIN DIA111
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3118.660 0.000 3119.780 1.120 ;
  LAYER metal4 ;
  RECT 3118.660 0.000 3119.780 1.120 ;
  LAYER metal3 ;
  RECT 3118.660 0.000 3119.780 1.120 ;
  LAYER metal2 ;
  RECT 3118.660 0.000 3119.780 1.120 ;
  LAYER metal1 ;
  RECT 3118.660 0.000 3119.780 1.120 ;
 END
END DIA111
PIN DOA111
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3105.640 0.000 3106.760 1.120 ;
  LAYER metal4 ;
  RECT 3105.640 0.000 3106.760 1.120 ;
  LAYER metal3 ;
  RECT 3105.640 0.000 3106.760 1.120 ;
  LAYER metal2 ;
  RECT 3105.640 0.000 3106.760 1.120 ;
  LAYER metal1 ;
  RECT 3105.640 0.000 3106.760 1.120 ;
 END
END DOA111
PIN DIA110
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3092.000 0.000 3093.120 1.120 ;
  LAYER metal4 ;
  RECT 3092.000 0.000 3093.120 1.120 ;
  LAYER metal3 ;
  RECT 3092.000 0.000 3093.120 1.120 ;
  LAYER metal2 ;
  RECT 3092.000 0.000 3093.120 1.120 ;
  LAYER metal1 ;
  RECT 3092.000 0.000 3093.120 1.120 ;
 END
END DIA110
PIN DOA110
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3078.360 0.000 3079.480 1.120 ;
  LAYER metal4 ;
  RECT 3078.360 0.000 3079.480 1.120 ;
  LAYER metal3 ;
  RECT 3078.360 0.000 3079.480 1.120 ;
  LAYER metal2 ;
  RECT 3078.360 0.000 3079.480 1.120 ;
  LAYER metal1 ;
  RECT 3078.360 0.000 3079.480 1.120 ;
 END
END DOA110
PIN DIA109
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 3065.340 0.000 3066.460 1.120 ;
  LAYER metal4 ;
  RECT 3065.340 0.000 3066.460 1.120 ;
  LAYER metal3 ;
  RECT 3065.340 0.000 3066.460 1.120 ;
  LAYER metal2 ;
  RECT 3065.340 0.000 3066.460 1.120 ;
  LAYER metal1 ;
  RECT 3065.340 0.000 3066.460 1.120 ;
 END
END DIA109
PIN DOA109
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 3051.700 0.000 3052.820 1.120 ;
  LAYER metal4 ;
  RECT 3051.700 0.000 3052.820 1.120 ;
  LAYER metal3 ;
  RECT 3051.700 0.000 3052.820 1.120 ;
  LAYER metal2 ;
  RECT 3051.700 0.000 3052.820 1.120 ;
  LAYER metal1 ;
  RECT 3051.700 0.000 3052.820 1.120 ;
 END
END DOA109
PIN DIA108
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3038.060 0.000 3039.180 1.120 ;
  LAYER metal4 ;
  RECT 3038.060 0.000 3039.180 1.120 ;
  LAYER metal3 ;
  RECT 3038.060 0.000 3039.180 1.120 ;
  LAYER metal2 ;
  RECT 3038.060 0.000 3039.180 1.120 ;
  LAYER metal1 ;
  RECT 3038.060 0.000 3039.180 1.120 ;
 END
END DIA108
PIN DOA108
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 3024.420 0.000 3025.540 1.120 ;
  LAYER metal4 ;
  RECT 3024.420 0.000 3025.540 1.120 ;
  LAYER metal3 ;
  RECT 3024.420 0.000 3025.540 1.120 ;
  LAYER metal2 ;
  RECT 3024.420 0.000 3025.540 1.120 ;
  LAYER metal1 ;
  RECT 3024.420 0.000 3025.540 1.120 ;
 END
END DOA108
PIN DIA107
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 3011.400 0.000 3012.520 1.120 ;
  LAYER metal4 ;
  RECT 3011.400 0.000 3012.520 1.120 ;
  LAYER metal3 ;
  RECT 3011.400 0.000 3012.520 1.120 ;
  LAYER metal2 ;
  RECT 3011.400 0.000 3012.520 1.120 ;
  LAYER metal1 ;
  RECT 3011.400 0.000 3012.520 1.120 ;
 END
END DIA107
PIN DOA107
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2997.760 0.000 2998.880 1.120 ;
  LAYER metal4 ;
  RECT 2997.760 0.000 2998.880 1.120 ;
  LAYER metal3 ;
  RECT 2997.760 0.000 2998.880 1.120 ;
  LAYER metal2 ;
  RECT 2997.760 0.000 2998.880 1.120 ;
  LAYER metal1 ;
  RECT 2997.760 0.000 2998.880 1.120 ;
 END
END DOA107
PIN DIA106
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2984.120 0.000 2985.240 1.120 ;
  LAYER metal4 ;
  RECT 2984.120 0.000 2985.240 1.120 ;
  LAYER metal3 ;
  RECT 2984.120 0.000 2985.240 1.120 ;
  LAYER metal2 ;
  RECT 2984.120 0.000 2985.240 1.120 ;
  LAYER metal1 ;
  RECT 2984.120 0.000 2985.240 1.120 ;
 END
END DIA106
PIN DOA106
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2971.100 0.000 2972.220 1.120 ;
  LAYER metal4 ;
  RECT 2971.100 0.000 2972.220 1.120 ;
  LAYER metal3 ;
  RECT 2971.100 0.000 2972.220 1.120 ;
  LAYER metal2 ;
  RECT 2971.100 0.000 2972.220 1.120 ;
  LAYER metal1 ;
  RECT 2971.100 0.000 2972.220 1.120 ;
 END
END DOA106
PIN DIA105
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2957.460 0.000 2958.580 1.120 ;
  LAYER metal4 ;
  RECT 2957.460 0.000 2958.580 1.120 ;
  LAYER metal3 ;
  RECT 2957.460 0.000 2958.580 1.120 ;
  LAYER metal2 ;
  RECT 2957.460 0.000 2958.580 1.120 ;
  LAYER metal1 ;
  RECT 2957.460 0.000 2958.580 1.120 ;
 END
END DIA105
PIN DOA105
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2943.820 0.000 2944.940 1.120 ;
  LAYER metal4 ;
  RECT 2943.820 0.000 2944.940 1.120 ;
  LAYER metal3 ;
  RECT 2943.820 0.000 2944.940 1.120 ;
  LAYER metal2 ;
  RECT 2943.820 0.000 2944.940 1.120 ;
  LAYER metal1 ;
  RECT 2943.820 0.000 2944.940 1.120 ;
 END
END DOA105
PIN DIA104
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2930.800 0.000 2931.920 1.120 ;
  LAYER metal4 ;
  RECT 2930.800 0.000 2931.920 1.120 ;
  LAYER metal3 ;
  RECT 2930.800 0.000 2931.920 1.120 ;
  LAYER metal2 ;
  RECT 2930.800 0.000 2931.920 1.120 ;
  LAYER metal1 ;
  RECT 2930.800 0.000 2931.920 1.120 ;
 END
END DIA104
PIN DOA104
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2917.160 0.000 2918.280 1.120 ;
  LAYER metal4 ;
  RECT 2917.160 0.000 2918.280 1.120 ;
  LAYER metal3 ;
  RECT 2917.160 0.000 2918.280 1.120 ;
  LAYER metal2 ;
  RECT 2917.160 0.000 2918.280 1.120 ;
  LAYER metal1 ;
  RECT 2917.160 0.000 2918.280 1.120 ;
 END
END DOA104
PIN DIA103
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2903.520 0.000 2904.640 1.120 ;
  LAYER metal4 ;
  RECT 2903.520 0.000 2904.640 1.120 ;
  LAYER metal3 ;
  RECT 2903.520 0.000 2904.640 1.120 ;
  LAYER metal2 ;
  RECT 2903.520 0.000 2904.640 1.120 ;
  LAYER metal1 ;
  RECT 2903.520 0.000 2904.640 1.120 ;
 END
END DIA103
PIN DOA103
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2890.500 0.000 2891.620 1.120 ;
  LAYER metal4 ;
  RECT 2890.500 0.000 2891.620 1.120 ;
  LAYER metal3 ;
  RECT 2890.500 0.000 2891.620 1.120 ;
  LAYER metal2 ;
  RECT 2890.500 0.000 2891.620 1.120 ;
  LAYER metal1 ;
  RECT 2890.500 0.000 2891.620 1.120 ;
 END
END DOA103
PIN DIA102
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2876.860 0.000 2877.980 1.120 ;
  LAYER metal4 ;
  RECT 2876.860 0.000 2877.980 1.120 ;
  LAYER metal3 ;
  RECT 2876.860 0.000 2877.980 1.120 ;
  LAYER metal2 ;
  RECT 2876.860 0.000 2877.980 1.120 ;
  LAYER metal1 ;
  RECT 2876.860 0.000 2877.980 1.120 ;
 END
END DIA102
PIN DOA102
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2863.220 0.000 2864.340 1.120 ;
  LAYER metal4 ;
  RECT 2863.220 0.000 2864.340 1.120 ;
  LAYER metal3 ;
  RECT 2863.220 0.000 2864.340 1.120 ;
  LAYER metal2 ;
  RECT 2863.220 0.000 2864.340 1.120 ;
  LAYER metal1 ;
  RECT 2863.220 0.000 2864.340 1.120 ;
 END
END DOA102
PIN DIA101
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2850.200 0.000 2851.320 1.120 ;
  LAYER metal4 ;
  RECT 2850.200 0.000 2851.320 1.120 ;
  LAYER metal3 ;
  RECT 2850.200 0.000 2851.320 1.120 ;
  LAYER metal2 ;
  RECT 2850.200 0.000 2851.320 1.120 ;
  LAYER metal1 ;
  RECT 2850.200 0.000 2851.320 1.120 ;
 END
END DIA101
PIN DOA101
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2836.560 0.000 2837.680 1.120 ;
  LAYER metal4 ;
  RECT 2836.560 0.000 2837.680 1.120 ;
  LAYER metal3 ;
  RECT 2836.560 0.000 2837.680 1.120 ;
  LAYER metal2 ;
  RECT 2836.560 0.000 2837.680 1.120 ;
  LAYER metal1 ;
  RECT 2836.560 0.000 2837.680 1.120 ;
 END
END DOA101
PIN DIA100
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2822.920 0.000 2824.040 1.120 ;
  LAYER metal4 ;
  RECT 2822.920 0.000 2824.040 1.120 ;
  LAYER metal3 ;
  RECT 2822.920 0.000 2824.040 1.120 ;
  LAYER metal2 ;
  RECT 2822.920 0.000 2824.040 1.120 ;
  LAYER metal1 ;
  RECT 2822.920 0.000 2824.040 1.120 ;
 END
END DIA100
PIN DOA100
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2809.900 0.000 2811.020 1.120 ;
  LAYER metal4 ;
  RECT 2809.900 0.000 2811.020 1.120 ;
  LAYER metal3 ;
  RECT 2809.900 0.000 2811.020 1.120 ;
  LAYER metal2 ;
  RECT 2809.900 0.000 2811.020 1.120 ;
  LAYER metal1 ;
  RECT 2809.900 0.000 2811.020 1.120 ;
 END
END DOA100
PIN DIA99
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2796.260 0.000 2797.380 1.120 ;
  LAYER metal4 ;
  RECT 2796.260 0.000 2797.380 1.120 ;
  LAYER metal3 ;
  RECT 2796.260 0.000 2797.380 1.120 ;
  LAYER metal2 ;
  RECT 2796.260 0.000 2797.380 1.120 ;
  LAYER metal1 ;
  RECT 2796.260 0.000 2797.380 1.120 ;
 END
END DIA99
PIN DOA99
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2782.620 0.000 2783.740 1.120 ;
  LAYER metal4 ;
  RECT 2782.620 0.000 2783.740 1.120 ;
  LAYER metal3 ;
  RECT 2782.620 0.000 2783.740 1.120 ;
  LAYER metal2 ;
  RECT 2782.620 0.000 2783.740 1.120 ;
  LAYER metal1 ;
  RECT 2782.620 0.000 2783.740 1.120 ;
 END
END DOA99
PIN DIA98
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2769.600 0.000 2770.720 1.120 ;
  LAYER metal4 ;
  RECT 2769.600 0.000 2770.720 1.120 ;
  LAYER metal3 ;
  RECT 2769.600 0.000 2770.720 1.120 ;
  LAYER metal2 ;
  RECT 2769.600 0.000 2770.720 1.120 ;
  LAYER metal1 ;
  RECT 2769.600 0.000 2770.720 1.120 ;
 END
END DIA98
PIN DOA98
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2755.960 0.000 2757.080 1.120 ;
  LAYER metal4 ;
  RECT 2755.960 0.000 2757.080 1.120 ;
  LAYER metal3 ;
  RECT 2755.960 0.000 2757.080 1.120 ;
  LAYER metal2 ;
  RECT 2755.960 0.000 2757.080 1.120 ;
  LAYER metal1 ;
  RECT 2755.960 0.000 2757.080 1.120 ;
 END
END DOA98
PIN DIA97
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2742.320 0.000 2743.440 1.120 ;
  LAYER metal4 ;
  RECT 2742.320 0.000 2743.440 1.120 ;
  LAYER metal3 ;
  RECT 2742.320 0.000 2743.440 1.120 ;
  LAYER metal2 ;
  RECT 2742.320 0.000 2743.440 1.120 ;
  LAYER metal1 ;
  RECT 2742.320 0.000 2743.440 1.120 ;
 END
END DIA97
PIN DOA97
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2729.300 0.000 2730.420 1.120 ;
  LAYER metal4 ;
  RECT 2729.300 0.000 2730.420 1.120 ;
  LAYER metal3 ;
  RECT 2729.300 0.000 2730.420 1.120 ;
  LAYER metal2 ;
  RECT 2729.300 0.000 2730.420 1.120 ;
  LAYER metal1 ;
  RECT 2729.300 0.000 2730.420 1.120 ;
 END
END DOA97
PIN DIA96
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2715.660 0.000 2716.780 1.120 ;
  LAYER metal4 ;
  RECT 2715.660 0.000 2716.780 1.120 ;
  LAYER metal3 ;
  RECT 2715.660 0.000 2716.780 1.120 ;
  LAYER metal2 ;
  RECT 2715.660 0.000 2716.780 1.120 ;
  LAYER metal1 ;
  RECT 2715.660 0.000 2716.780 1.120 ;
 END
END DIA96
PIN DOA96
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2702.020 0.000 2703.140 1.120 ;
  LAYER metal4 ;
  RECT 2702.020 0.000 2703.140 1.120 ;
  LAYER metal3 ;
  RECT 2702.020 0.000 2703.140 1.120 ;
  LAYER metal2 ;
  RECT 2702.020 0.000 2703.140 1.120 ;
  LAYER metal1 ;
  RECT 2702.020 0.000 2703.140 1.120 ;
 END
END DOA96
PIN DIA95
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2689.000 0.000 2690.120 1.120 ;
  LAYER metal4 ;
  RECT 2689.000 0.000 2690.120 1.120 ;
  LAYER metal3 ;
  RECT 2689.000 0.000 2690.120 1.120 ;
  LAYER metal2 ;
  RECT 2689.000 0.000 2690.120 1.120 ;
  LAYER metal1 ;
  RECT 2689.000 0.000 2690.120 1.120 ;
 END
END DIA95
PIN DOA95
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2675.360 0.000 2676.480 1.120 ;
  LAYER metal4 ;
  RECT 2675.360 0.000 2676.480 1.120 ;
  LAYER metal3 ;
  RECT 2675.360 0.000 2676.480 1.120 ;
  LAYER metal2 ;
  RECT 2675.360 0.000 2676.480 1.120 ;
  LAYER metal1 ;
  RECT 2675.360 0.000 2676.480 1.120 ;
 END
END DOA95
PIN DIA94
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2661.720 0.000 2662.840 1.120 ;
  LAYER metal4 ;
  RECT 2661.720 0.000 2662.840 1.120 ;
  LAYER metal3 ;
  RECT 2661.720 0.000 2662.840 1.120 ;
  LAYER metal2 ;
  RECT 2661.720 0.000 2662.840 1.120 ;
  LAYER metal1 ;
  RECT 2661.720 0.000 2662.840 1.120 ;
 END
END DIA94
PIN DOA94
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2648.700 0.000 2649.820 1.120 ;
  LAYER metal4 ;
  RECT 2648.700 0.000 2649.820 1.120 ;
  LAYER metal3 ;
  RECT 2648.700 0.000 2649.820 1.120 ;
  LAYER metal2 ;
  RECT 2648.700 0.000 2649.820 1.120 ;
  LAYER metal1 ;
  RECT 2648.700 0.000 2649.820 1.120 ;
 END
END DOA94
PIN DIA93
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2635.060 0.000 2636.180 1.120 ;
  LAYER metal4 ;
  RECT 2635.060 0.000 2636.180 1.120 ;
  LAYER metal3 ;
  RECT 2635.060 0.000 2636.180 1.120 ;
  LAYER metal2 ;
  RECT 2635.060 0.000 2636.180 1.120 ;
  LAYER metal1 ;
  RECT 2635.060 0.000 2636.180 1.120 ;
 END
END DIA93
PIN DOA93
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2621.420 0.000 2622.540 1.120 ;
  LAYER metal4 ;
  RECT 2621.420 0.000 2622.540 1.120 ;
  LAYER metal3 ;
  RECT 2621.420 0.000 2622.540 1.120 ;
  LAYER metal2 ;
  RECT 2621.420 0.000 2622.540 1.120 ;
  LAYER metal1 ;
  RECT 2621.420 0.000 2622.540 1.120 ;
 END
END DOA93
PIN DIA92
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2607.780 0.000 2608.900 1.120 ;
  LAYER metal4 ;
  RECT 2607.780 0.000 2608.900 1.120 ;
  LAYER metal3 ;
  RECT 2607.780 0.000 2608.900 1.120 ;
  LAYER metal2 ;
  RECT 2607.780 0.000 2608.900 1.120 ;
  LAYER metal1 ;
  RECT 2607.780 0.000 2608.900 1.120 ;
 END
END DIA92
PIN DOA92
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2594.760 0.000 2595.880 1.120 ;
  LAYER metal4 ;
  RECT 2594.760 0.000 2595.880 1.120 ;
  LAYER metal3 ;
  RECT 2594.760 0.000 2595.880 1.120 ;
  LAYER metal2 ;
  RECT 2594.760 0.000 2595.880 1.120 ;
  LAYER metal1 ;
  RECT 2594.760 0.000 2595.880 1.120 ;
 END
END DOA92
PIN DIA91
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2581.120 0.000 2582.240 1.120 ;
  LAYER metal4 ;
  RECT 2581.120 0.000 2582.240 1.120 ;
  LAYER metal3 ;
  RECT 2581.120 0.000 2582.240 1.120 ;
  LAYER metal2 ;
  RECT 2581.120 0.000 2582.240 1.120 ;
  LAYER metal1 ;
  RECT 2581.120 0.000 2582.240 1.120 ;
 END
END DIA91
PIN DOA91
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2567.480 0.000 2568.600 1.120 ;
  LAYER metal4 ;
  RECT 2567.480 0.000 2568.600 1.120 ;
  LAYER metal3 ;
  RECT 2567.480 0.000 2568.600 1.120 ;
  LAYER metal2 ;
  RECT 2567.480 0.000 2568.600 1.120 ;
  LAYER metal1 ;
  RECT 2567.480 0.000 2568.600 1.120 ;
 END
END DOA91
PIN DIA90
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2554.460 0.000 2555.580 1.120 ;
  LAYER metal4 ;
  RECT 2554.460 0.000 2555.580 1.120 ;
  LAYER metal3 ;
  RECT 2554.460 0.000 2555.580 1.120 ;
  LAYER metal2 ;
  RECT 2554.460 0.000 2555.580 1.120 ;
  LAYER metal1 ;
  RECT 2554.460 0.000 2555.580 1.120 ;
 END
END DIA90
PIN DOA90
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2540.820 0.000 2541.940 1.120 ;
  LAYER metal4 ;
  RECT 2540.820 0.000 2541.940 1.120 ;
  LAYER metal3 ;
  RECT 2540.820 0.000 2541.940 1.120 ;
  LAYER metal2 ;
  RECT 2540.820 0.000 2541.940 1.120 ;
  LAYER metal1 ;
  RECT 2540.820 0.000 2541.940 1.120 ;
 END
END DOA90
PIN DIA89
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2527.180 0.000 2528.300 1.120 ;
  LAYER metal4 ;
  RECT 2527.180 0.000 2528.300 1.120 ;
  LAYER metal3 ;
  RECT 2527.180 0.000 2528.300 1.120 ;
  LAYER metal2 ;
  RECT 2527.180 0.000 2528.300 1.120 ;
  LAYER metal1 ;
  RECT 2527.180 0.000 2528.300 1.120 ;
 END
END DIA89
PIN DOA89
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2514.160 0.000 2515.280 1.120 ;
  LAYER metal4 ;
  RECT 2514.160 0.000 2515.280 1.120 ;
  LAYER metal3 ;
  RECT 2514.160 0.000 2515.280 1.120 ;
  LAYER metal2 ;
  RECT 2514.160 0.000 2515.280 1.120 ;
  LAYER metal1 ;
  RECT 2514.160 0.000 2515.280 1.120 ;
 END
END DOA89
PIN DIA88
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2500.520 0.000 2501.640 1.120 ;
  LAYER metal4 ;
  RECT 2500.520 0.000 2501.640 1.120 ;
  LAYER metal3 ;
  RECT 2500.520 0.000 2501.640 1.120 ;
  LAYER metal2 ;
  RECT 2500.520 0.000 2501.640 1.120 ;
  LAYER metal1 ;
  RECT 2500.520 0.000 2501.640 1.120 ;
 END
END DIA88
PIN DOA88
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2486.880 0.000 2488.000 1.120 ;
  LAYER metal4 ;
  RECT 2486.880 0.000 2488.000 1.120 ;
  LAYER metal3 ;
  RECT 2486.880 0.000 2488.000 1.120 ;
  LAYER metal2 ;
  RECT 2486.880 0.000 2488.000 1.120 ;
  LAYER metal1 ;
  RECT 2486.880 0.000 2488.000 1.120 ;
 END
END DOA88
PIN DIA87
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2473.860 0.000 2474.980 1.120 ;
  LAYER metal4 ;
  RECT 2473.860 0.000 2474.980 1.120 ;
  LAYER metal3 ;
  RECT 2473.860 0.000 2474.980 1.120 ;
  LAYER metal2 ;
  RECT 2473.860 0.000 2474.980 1.120 ;
  LAYER metal1 ;
  RECT 2473.860 0.000 2474.980 1.120 ;
 END
END DIA87
PIN DOA87
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2460.220 0.000 2461.340 1.120 ;
  LAYER metal4 ;
  RECT 2460.220 0.000 2461.340 1.120 ;
  LAYER metal3 ;
  RECT 2460.220 0.000 2461.340 1.120 ;
  LAYER metal2 ;
  RECT 2460.220 0.000 2461.340 1.120 ;
  LAYER metal1 ;
  RECT 2460.220 0.000 2461.340 1.120 ;
 END
END DOA87
PIN DIA86
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2446.580 0.000 2447.700 1.120 ;
  LAYER metal4 ;
  RECT 2446.580 0.000 2447.700 1.120 ;
  LAYER metal3 ;
  RECT 2446.580 0.000 2447.700 1.120 ;
  LAYER metal2 ;
  RECT 2446.580 0.000 2447.700 1.120 ;
  LAYER metal1 ;
  RECT 2446.580 0.000 2447.700 1.120 ;
 END
END DIA86
PIN DOA86
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2433.560 0.000 2434.680 1.120 ;
  LAYER metal4 ;
  RECT 2433.560 0.000 2434.680 1.120 ;
  LAYER metal3 ;
  RECT 2433.560 0.000 2434.680 1.120 ;
  LAYER metal2 ;
  RECT 2433.560 0.000 2434.680 1.120 ;
  LAYER metal1 ;
  RECT 2433.560 0.000 2434.680 1.120 ;
 END
END DOA86
PIN DIA85
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2419.920 0.000 2421.040 1.120 ;
  LAYER metal4 ;
  RECT 2419.920 0.000 2421.040 1.120 ;
  LAYER metal3 ;
  RECT 2419.920 0.000 2421.040 1.120 ;
  LAYER metal2 ;
  RECT 2419.920 0.000 2421.040 1.120 ;
  LAYER metal1 ;
  RECT 2419.920 0.000 2421.040 1.120 ;
 END
END DIA85
PIN DOA85
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2406.280 0.000 2407.400 1.120 ;
  LAYER metal4 ;
  RECT 2406.280 0.000 2407.400 1.120 ;
  LAYER metal3 ;
  RECT 2406.280 0.000 2407.400 1.120 ;
  LAYER metal2 ;
  RECT 2406.280 0.000 2407.400 1.120 ;
  LAYER metal1 ;
  RECT 2406.280 0.000 2407.400 1.120 ;
 END
END DOA85
PIN DIA84
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2393.260 0.000 2394.380 1.120 ;
  LAYER metal4 ;
  RECT 2393.260 0.000 2394.380 1.120 ;
  LAYER metal3 ;
  RECT 2393.260 0.000 2394.380 1.120 ;
  LAYER metal2 ;
  RECT 2393.260 0.000 2394.380 1.120 ;
  LAYER metal1 ;
  RECT 2393.260 0.000 2394.380 1.120 ;
 END
END DIA84
PIN DOA84
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2379.620 0.000 2380.740 1.120 ;
  LAYER metal4 ;
  RECT 2379.620 0.000 2380.740 1.120 ;
  LAYER metal3 ;
  RECT 2379.620 0.000 2380.740 1.120 ;
  LAYER metal2 ;
  RECT 2379.620 0.000 2380.740 1.120 ;
  LAYER metal1 ;
  RECT 2379.620 0.000 2380.740 1.120 ;
 END
END DOA84
PIN DIA83
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2365.980 0.000 2367.100 1.120 ;
  LAYER metal4 ;
  RECT 2365.980 0.000 2367.100 1.120 ;
  LAYER metal3 ;
  RECT 2365.980 0.000 2367.100 1.120 ;
  LAYER metal2 ;
  RECT 2365.980 0.000 2367.100 1.120 ;
  LAYER metal1 ;
  RECT 2365.980 0.000 2367.100 1.120 ;
 END
END DIA83
PIN DOA83
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2352.960 0.000 2354.080 1.120 ;
  LAYER metal4 ;
  RECT 2352.960 0.000 2354.080 1.120 ;
  LAYER metal3 ;
  RECT 2352.960 0.000 2354.080 1.120 ;
  LAYER metal2 ;
  RECT 2352.960 0.000 2354.080 1.120 ;
  LAYER metal1 ;
  RECT 2352.960 0.000 2354.080 1.120 ;
 END
END DOA83
PIN DIA82
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2339.320 0.000 2340.440 1.120 ;
  LAYER metal4 ;
  RECT 2339.320 0.000 2340.440 1.120 ;
  LAYER metal3 ;
  RECT 2339.320 0.000 2340.440 1.120 ;
  LAYER metal2 ;
  RECT 2339.320 0.000 2340.440 1.120 ;
  LAYER metal1 ;
  RECT 2339.320 0.000 2340.440 1.120 ;
 END
END DIA82
PIN DOA82
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2325.680 0.000 2326.800 1.120 ;
  LAYER metal4 ;
  RECT 2325.680 0.000 2326.800 1.120 ;
  LAYER metal3 ;
  RECT 2325.680 0.000 2326.800 1.120 ;
  LAYER metal2 ;
  RECT 2325.680 0.000 2326.800 1.120 ;
  LAYER metal1 ;
  RECT 2325.680 0.000 2326.800 1.120 ;
 END
END DOA82
PIN DIA81
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2312.660 0.000 2313.780 1.120 ;
  LAYER metal4 ;
  RECT 2312.660 0.000 2313.780 1.120 ;
  LAYER metal3 ;
  RECT 2312.660 0.000 2313.780 1.120 ;
  LAYER metal2 ;
  RECT 2312.660 0.000 2313.780 1.120 ;
  LAYER metal1 ;
  RECT 2312.660 0.000 2313.780 1.120 ;
 END
END DIA81
PIN DOA81
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2299.020 0.000 2300.140 1.120 ;
  LAYER metal4 ;
  RECT 2299.020 0.000 2300.140 1.120 ;
  LAYER metal3 ;
  RECT 2299.020 0.000 2300.140 1.120 ;
  LAYER metal2 ;
  RECT 2299.020 0.000 2300.140 1.120 ;
  LAYER metal1 ;
  RECT 2299.020 0.000 2300.140 1.120 ;
 END
END DOA81
PIN DIA80
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2285.380 0.000 2286.500 1.120 ;
  LAYER metal4 ;
  RECT 2285.380 0.000 2286.500 1.120 ;
  LAYER metal3 ;
  RECT 2285.380 0.000 2286.500 1.120 ;
  LAYER metal2 ;
  RECT 2285.380 0.000 2286.500 1.120 ;
  LAYER metal1 ;
  RECT 2285.380 0.000 2286.500 1.120 ;
 END
END DIA80
PIN DOA80
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2272.360 0.000 2273.480 1.120 ;
  LAYER metal4 ;
  RECT 2272.360 0.000 2273.480 1.120 ;
  LAYER metal3 ;
  RECT 2272.360 0.000 2273.480 1.120 ;
  LAYER metal2 ;
  RECT 2272.360 0.000 2273.480 1.120 ;
  LAYER metal1 ;
  RECT 2272.360 0.000 2273.480 1.120 ;
 END
END DOA80
PIN DIA79
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2258.720 0.000 2259.840 1.120 ;
  LAYER metal4 ;
  RECT 2258.720 0.000 2259.840 1.120 ;
  LAYER metal3 ;
  RECT 2258.720 0.000 2259.840 1.120 ;
  LAYER metal2 ;
  RECT 2258.720 0.000 2259.840 1.120 ;
  LAYER metal1 ;
  RECT 2258.720 0.000 2259.840 1.120 ;
 END
END DIA79
PIN DOA79
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2245.080 0.000 2246.200 1.120 ;
  LAYER metal4 ;
  RECT 2245.080 0.000 2246.200 1.120 ;
  LAYER metal3 ;
  RECT 2245.080 0.000 2246.200 1.120 ;
  LAYER metal2 ;
  RECT 2245.080 0.000 2246.200 1.120 ;
  LAYER metal1 ;
  RECT 2245.080 0.000 2246.200 1.120 ;
 END
END DOA79
PIN DIA78
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2232.060 0.000 2233.180 1.120 ;
  LAYER metal4 ;
  RECT 2232.060 0.000 2233.180 1.120 ;
  LAYER metal3 ;
  RECT 2232.060 0.000 2233.180 1.120 ;
  LAYER metal2 ;
  RECT 2232.060 0.000 2233.180 1.120 ;
  LAYER metal1 ;
  RECT 2232.060 0.000 2233.180 1.120 ;
 END
END DIA78
PIN DOA78
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2218.420 0.000 2219.540 1.120 ;
  LAYER metal4 ;
  RECT 2218.420 0.000 2219.540 1.120 ;
  LAYER metal3 ;
  RECT 2218.420 0.000 2219.540 1.120 ;
  LAYER metal2 ;
  RECT 2218.420 0.000 2219.540 1.120 ;
  LAYER metal1 ;
  RECT 2218.420 0.000 2219.540 1.120 ;
 END
END DOA78
PIN DIA77
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2204.780 0.000 2205.900 1.120 ;
  LAYER metal4 ;
  RECT 2204.780 0.000 2205.900 1.120 ;
  LAYER metal3 ;
  RECT 2204.780 0.000 2205.900 1.120 ;
  LAYER metal2 ;
  RECT 2204.780 0.000 2205.900 1.120 ;
  LAYER metal1 ;
  RECT 2204.780 0.000 2205.900 1.120 ;
 END
END DIA77
PIN DOA77
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2191.140 0.000 2192.260 1.120 ;
  LAYER metal4 ;
  RECT 2191.140 0.000 2192.260 1.120 ;
  LAYER metal3 ;
  RECT 2191.140 0.000 2192.260 1.120 ;
  LAYER metal2 ;
  RECT 2191.140 0.000 2192.260 1.120 ;
  LAYER metal1 ;
  RECT 2191.140 0.000 2192.260 1.120 ;
 END
END DOA77
PIN DIA76
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2178.120 0.000 2179.240 1.120 ;
  LAYER metal4 ;
  RECT 2178.120 0.000 2179.240 1.120 ;
  LAYER metal3 ;
  RECT 2178.120 0.000 2179.240 1.120 ;
  LAYER metal2 ;
  RECT 2178.120 0.000 2179.240 1.120 ;
  LAYER metal1 ;
  RECT 2178.120 0.000 2179.240 1.120 ;
 END
END DIA76
PIN DOA76
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2164.480 0.000 2165.600 1.120 ;
  LAYER metal4 ;
  RECT 2164.480 0.000 2165.600 1.120 ;
  LAYER metal3 ;
  RECT 2164.480 0.000 2165.600 1.120 ;
  LAYER metal2 ;
  RECT 2164.480 0.000 2165.600 1.120 ;
  LAYER metal1 ;
  RECT 2164.480 0.000 2165.600 1.120 ;
 END
END DOA76
PIN DIA75
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2150.840 0.000 2151.960 1.120 ;
  LAYER metal4 ;
  RECT 2150.840 0.000 2151.960 1.120 ;
  LAYER metal3 ;
  RECT 2150.840 0.000 2151.960 1.120 ;
  LAYER metal2 ;
  RECT 2150.840 0.000 2151.960 1.120 ;
  LAYER metal1 ;
  RECT 2150.840 0.000 2151.960 1.120 ;
 END
END DIA75
PIN DOA75
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2137.820 0.000 2138.940 1.120 ;
  LAYER metal4 ;
  RECT 2137.820 0.000 2138.940 1.120 ;
  LAYER metal3 ;
  RECT 2137.820 0.000 2138.940 1.120 ;
  LAYER metal2 ;
  RECT 2137.820 0.000 2138.940 1.120 ;
  LAYER metal1 ;
  RECT 2137.820 0.000 2138.940 1.120 ;
 END
END DOA75
PIN DIA74
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2124.180 0.000 2125.300 1.120 ;
  LAYER metal4 ;
  RECT 2124.180 0.000 2125.300 1.120 ;
  LAYER metal3 ;
  RECT 2124.180 0.000 2125.300 1.120 ;
  LAYER metal2 ;
  RECT 2124.180 0.000 2125.300 1.120 ;
  LAYER metal1 ;
  RECT 2124.180 0.000 2125.300 1.120 ;
 END
END DIA74
PIN DOA74
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2110.540 0.000 2111.660 1.120 ;
  LAYER metal4 ;
  RECT 2110.540 0.000 2111.660 1.120 ;
  LAYER metal3 ;
  RECT 2110.540 0.000 2111.660 1.120 ;
  LAYER metal2 ;
  RECT 2110.540 0.000 2111.660 1.120 ;
  LAYER metal1 ;
  RECT 2110.540 0.000 2111.660 1.120 ;
 END
END DOA74
PIN DIA73
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2097.520 0.000 2098.640 1.120 ;
  LAYER metal4 ;
  RECT 2097.520 0.000 2098.640 1.120 ;
  LAYER metal3 ;
  RECT 2097.520 0.000 2098.640 1.120 ;
  LAYER metal2 ;
  RECT 2097.520 0.000 2098.640 1.120 ;
  LAYER metal1 ;
  RECT 2097.520 0.000 2098.640 1.120 ;
 END
END DIA73
PIN DOA73
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2083.880 0.000 2085.000 1.120 ;
  LAYER metal4 ;
  RECT 2083.880 0.000 2085.000 1.120 ;
  LAYER metal3 ;
  RECT 2083.880 0.000 2085.000 1.120 ;
  LAYER metal2 ;
  RECT 2083.880 0.000 2085.000 1.120 ;
  LAYER metal1 ;
  RECT 2083.880 0.000 2085.000 1.120 ;
 END
END DOA73
PIN DIA72
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2070.240 0.000 2071.360 1.120 ;
  LAYER metal4 ;
  RECT 2070.240 0.000 2071.360 1.120 ;
  LAYER metal3 ;
  RECT 2070.240 0.000 2071.360 1.120 ;
  LAYER metal2 ;
  RECT 2070.240 0.000 2071.360 1.120 ;
  LAYER metal1 ;
  RECT 2070.240 0.000 2071.360 1.120 ;
 END
END DIA72
PIN DOA72
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2057.220 0.000 2058.340 1.120 ;
  LAYER metal4 ;
  RECT 2057.220 0.000 2058.340 1.120 ;
  LAYER metal3 ;
  RECT 2057.220 0.000 2058.340 1.120 ;
  LAYER metal2 ;
  RECT 2057.220 0.000 2058.340 1.120 ;
  LAYER metal1 ;
  RECT 2057.220 0.000 2058.340 1.120 ;
 END
END DOA72
PIN DIA71
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 2043.580 0.000 2044.700 1.120 ;
  LAYER metal4 ;
  RECT 2043.580 0.000 2044.700 1.120 ;
  LAYER metal3 ;
  RECT 2043.580 0.000 2044.700 1.120 ;
  LAYER metal2 ;
  RECT 2043.580 0.000 2044.700 1.120 ;
  LAYER metal1 ;
  RECT 2043.580 0.000 2044.700 1.120 ;
 END
END DIA71
PIN DOA71
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 2029.940 0.000 2031.060 1.120 ;
  LAYER metal4 ;
  RECT 2029.940 0.000 2031.060 1.120 ;
  LAYER metal3 ;
  RECT 2029.940 0.000 2031.060 1.120 ;
  LAYER metal2 ;
  RECT 2029.940 0.000 2031.060 1.120 ;
  LAYER metal1 ;
  RECT 2029.940 0.000 2031.060 1.120 ;
 END
END DOA71
PIN DIA70
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 2016.920 0.000 2018.040 1.120 ;
  LAYER metal4 ;
  RECT 2016.920 0.000 2018.040 1.120 ;
  LAYER metal3 ;
  RECT 2016.920 0.000 2018.040 1.120 ;
  LAYER metal2 ;
  RECT 2016.920 0.000 2018.040 1.120 ;
  LAYER metal1 ;
  RECT 2016.920 0.000 2018.040 1.120 ;
 END
END DIA70
PIN DOA70
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 2003.280 0.000 2004.400 1.120 ;
  LAYER metal4 ;
  RECT 2003.280 0.000 2004.400 1.120 ;
  LAYER metal3 ;
  RECT 2003.280 0.000 2004.400 1.120 ;
  LAYER metal2 ;
  RECT 2003.280 0.000 2004.400 1.120 ;
  LAYER metal1 ;
  RECT 2003.280 0.000 2004.400 1.120 ;
 END
END DOA70
PIN DIA69
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1989.640 0.000 1990.760 1.120 ;
  LAYER metal4 ;
  RECT 1989.640 0.000 1990.760 1.120 ;
  LAYER metal3 ;
  RECT 1989.640 0.000 1990.760 1.120 ;
  LAYER metal2 ;
  RECT 1989.640 0.000 1990.760 1.120 ;
  LAYER metal1 ;
  RECT 1989.640 0.000 1990.760 1.120 ;
 END
END DIA69
PIN DOA69
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1976.620 0.000 1977.740 1.120 ;
  LAYER metal4 ;
  RECT 1976.620 0.000 1977.740 1.120 ;
  LAYER metal3 ;
  RECT 1976.620 0.000 1977.740 1.120 ;
  LAYER metal2 ;
  RECT 1976.620 0.000 1977.740 1.120 ;
  LAYER metal1 ;
  RECT 1976.620 0.000 1977.740 1.120 ;
 END
END DOA69
PIN DIA68
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1962.980 0.000 1964.100 1.120 ;
  LAYER metal4 ;
  RECT 1962.980 0.000 1964.100 1.120 ;
  LAYER metal3 ;
  RECT 1962.980 0.000 1964.100 1.120 ;
  LAYER metal2 ;
  RECT 1962.980 0.000 1964.100 1.120 ;
  LAYER metal1 ;
  RECT 1962.980 0.000 1964.100 1.120 ;
 END
END DIA68
PIN DOA68
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1949.340 0.000 1950.460 1.120 ;
  LAYER metal4 ;
  RECT 1949.340 0.000 1950.460 1.120 ;
  LAYER metal3 ;
  RECT 1949.340 0.000 1950.460 1.120 ;
  LAYER metal2 ;
  RECT 1949.340 0.000 1950.460 1.120 ;
  LAYER metal1 ;
  RECT 1949.340 0.000 1950.460 1.120 ;
 END
END DOA68
PIN DIA67
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1936.320 0.000 1937.440 1.120 ;
  LAYER metal4 ;
  RECT 1936.320 0.000 1937.440 1.120 ;
  LAYER metal3 ;
  RECT 1936.320 0.000 1937.440 1.120 ;
  LAYER metal2 ;
  RECT 1936.320 0.000 1937.440 1.120 ;
  LAYER metal1 ;
  RECT 1936.320 0.000 1937.440 1.120 ;
 END
END DIA67
PIN DOA67
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1922.680 0.000 1923.800 1.120 ;
  LAYER metal4 ;
  RECT 1922.680 0.000 1923.800 1.120 ;
  LAYER metal3 ;
  RECT 1922.680 0.000 1923.800 1.120 ;
  LAYER metal2 ;
  RECT 1922.680 0.000 1923.800 1.120 ;
  LAYER metal1 ;
  RECT 1922.680 0.000 1923.800 1.120 ;
 END
END DOA67
PIN DIA66
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1909.040 0.000 1910.160 1.120 ;
  LAYER metal4 ;
  RECT 1909.040 0.000 1910.160 1.120 ;
  LAYER metal3 ;
  RECT 1909.040 0.000 1910.160 1.120 ;
  LAYER metal2 ;
  RECT 1909.040 0.000 1910.160 1.120 ;
  LAYER metal1 ;
  RECT 1909.040 0.000 1910.160 1.120 ;
 END
END DIA66
PIN DOA66
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1896.020 0.000 1897.140 1.120 ;
  LAYER metal4 ;
  RECT 1896.020 0.000 1897.140 1.120 ;
  LAYER metal3 ;
  RECT 1896.020 0.000 1897.140 1.120 ;
  LAYER metal2 ;
  RECT 1896.020 0.000 1897.140 1.120 ;
  LAYER metal1 ;
  RECT 1896.020 0.000 1897.140 1.120 ;
 END
END DOA66
PIN DIA65
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1882.380 0.000 1883.500 1.120 ;
  LAYER metal4 ;
  RECT 1882.380 0.000 1883.500 1.120 ;
  LAYER metal3 ;
  RECT 1882.380 0.000 1883.500 1.120 ;
  LAYER metal2 ;
  RECT 1882.380 0.000 1883.500 1.120 ;
  LAYER metal1 ;
  RECT 1882.380 0.000 1883.500 1.120 ;
 END
END DIA65
PIN DOA65
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1868.740 0.000 1869.860 1.120 ;
  LAYER metal4 ;
  RECT 1868.740 0.000 1869.860 1.120 ;
  LAYER metal3 ;
  RECT 1868.740 0.000 1869.860 1.120 ;
  LAYER metal2 ;
  RECT 1868.740 0.000 1869.860 1.120 ;
  LAYER metal1 ;
  RECT 1868.740 0.000 1869.860 1.120 ;
 END
END DOA65
PIN DIA64
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1855.720 0.000 1856.840 1.120 ;
  LAYER metal4 ;
  RECT 1855.720 0.000 1856.840 1.120 ;
  LAYER metal3 ;
  RECT 1855.720 0.000 1856.840 1.120 ;
  LAYER metal2 ;
  RECT 1855.720 0.000 1856.840 1.120 ;
  LAYER metal1 ;
  RECT 1855.720 0.000 1856.840 1.120 ;
 END
END DIA64
PIN DOA64
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1842.080 0.000 1843.200 1.120 ;
  LAYER metal4 ;
  RECT 1842.080 0.000 1843.200 1.120 ;
  LAYER metal3 ;
  RECT 1842.080 0.000 1843.200 1.120 ;
  LAYER metal2 ;
  RECT 1842.080 0.000 1843.200 1.120 ;
  LAYER metal1 ;
  RECT 1842.080 0.000 1843.200 1.120 ;
 END
END DOA64
PIN OEA
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1815.420 0.000 1816.540 1.120 ;
  LAYER metal4 ;
  RECT 1815.420 0.000 1816.540 1.120 ;
  LAYER metal3 ;
  RECT 1815.420 0.000 1816.540 1.120 ;
  LAYER metal2 ;
  RECT 1815.420 0.000 1816.540 1.120 ;
  LAYER metal1 ;
  RECT 1815.420 0.000 1816.540 1.120 ;
 END
END OEA
PIN CKA
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1801.780 0.000 1802.900 1.120 ;
  LAYER metal4 ;
  RECT 1801.780 0.000 1802.900 1.120 ;
  LAYER metal3 ;
  RECT 1801.780 0.000 1802.900 1.120 ;
  LAYER metal2 ;
  RECT 1801.780 0.000 1802.900 1.120 ;
  LAYER metal1 ;
  RECT 1801.780 0.000 1802.900 1.120 ;
 END
END CKA
PIN CSA
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1799.920 0.000 1801.040 1.120 ;
  LAYER metal4 ;
  RECT 1799.920 0.000 1801.040 1.120 ;
  LAYER metal3 ;
  RECT 1799.920 0.000 1801.040 1.120 ;
  LAYER metal2 ;
  RECT 1799.920 0.000 1801.040 1.120 ;
  LAYER metal1 ;
  RECT 1799.920 0.000 1801.040 1.120 ;
 END
END CSA
PIN WEAN
  DIRECTION INPUT ;
  CAPACITANCE 0.013 ;
 PORT
  LAYER metal5 ;
  RECT 1797.440 0.000 1798.560 1.120 ;
  LAYER metal4 ;
  RECT 1797.440 0.000 1798.560 1.120 ;
  LAYER metal3 ;
  RECT 1797.440 0.000 1798.560 1.120 ;
  LAYER metal2 ;
  RECT 1797.440 0.000 1798.560 1.120 ;
  LAYER metal1 ;
  RECT 1797.440 0.000 1798.560 1.120 ;
 END
END WEAN
PIN A2
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1793.720 0.000 1794.840 1.120 ;
  LAYER metal4 ;
  RECT 1793.720 0.000 1794.840 1.120 ;
  LAYER metal3 ;
  RECT 1793.720 0.000 1794.840 1.120 ;
  LAYER metal2 ;
  RECT 1793.720 0.000 1794.840 1.120 ;
  LAYER metal1 ;
  RECT 1793.720 0.000 1794.840 1.120 ;
 END
END A2
PIN A1
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1788.140 0.000 1789.260 1.120 ;
  LAYER metal4 ;
  RECT 1788.140 0.000 1789.260 1.120 ;
  LAYER metal3 ;
  RECT 1788.140 0.000 1789.260 1.120 ;
  LAYER metal2 ;
  RECT 1788.140 0.000 1789.260 1.120 ;
  LAYER metal1 ;
  RECT 1788.140 0.000 1789.260 1.120 ;
 END
END A1
PIN A0
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1786.280 0.000 1787.400 1.120 ;
  LAYER metal4 ;
  RECT 1786.280 0.000 1787.400 1.120 ;
  LAYER metal3 ;
  RECT 1786.280 0.000 1787.400 1.120 ;
  LAYER metal2 ;
  RECT 1786.280 0.000 1787.400 1.120 ;
  LAYER metal1 ;
  RECT 1786.280 0.000 1787.400 1.120 ;
 END
END A0
PIN A5
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1777.600 0.000 1778.720 1.120 ;
  LAYER metal4 ;
  RECT 1777.600 0.000 1778.720 1.120 ;
  LAYER metal3 ;
  RECT 1777.600 0.000 1778.720 1.120 ;
  LAYER metal2 ;
  RECT 1777.600 0.000 1778.720 1.120 ;
  LAYER metal1 ;
  RECT 1777.600 0.000 1778.720 1.120 ;
 END
END A5
PIN A4
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1772.020 0.000 1773.140 1.120 ;
  LAYER metal4 ;
  RECT 1772.020 0.000 1773.140 1.120 ;
  LAYER metal3 ;
  RECT 1772.020 0.000 1773.140 1.120 ;
  LAYER metal2 ;
  RECT 1772.020 0.000 1773.140 1.120 ;
  LAYER metal1 ;
  RECT 1772.020 0.000 1773.140 1.120 ;
 END
END A4
PIN A3
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1766.440 0.000 1767.560 1.120 ;
  LAYER metal4 ;
  RECT 1766.440 0.000 1767.560 1.120 ;
  LAYER metal3 ;
  RECT 1766.440 0.000 1767.560 1.120 ;
  LAYER metal2 ;
  RECT 1766.440 0.000 1767.560 1.120 ;
  LAYER metal1 ;
  RECT 1766.440 0.000 1767.560 1.120 ;
 END
END A3
PIN A7
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1747.840 0.000 1748.960 1.120 ;
  LAYER metal4 ;
  RECT 1747.840 0.000 1748.960 1.120 ;
  LAYER metal3 ;
  RECT 1747.840 0.000 1748.960 1.120 ;
  LAYER metal2 ;
  RECT 1747.840 0.000 1748.960 1.120 ;
  LAYER metal1 ;
  RECT 1747.840 0.000 1748.960 1.120 ;
 END
END A7
PIN A6
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1741.640 0.000 1742.760 1.120 ;
  LAYER metal4 ;
  RECT 1741.640 0.000 1742.760 1.120 ;
  LAYER metal3 ;
  RECT 1741.640 0.000 1742.760 1.120 ;
  LAYER metal2 ;
  RECT 1741.640 0.000 1742.760 1.120 ;
  LAYER metal1 ;
  RECT 1741.640 0.000 1742.760 1.120 ;
 END
END A6
PIN DIA63
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1719.320 0.000 1720.440 1.120 ;
  LAYER metal4 ;
  RECT 1719.320 0.000 1720.440 1.120 ;
  LAYER metal3 ;
  RECT 1719.320 0.000 1720.440 1.120 ;
  LAYER metal2 ;
  RECT 1719.320 0.000 1720.440 1.120 ;
  LAYER metal1 ;
  RECT 1719.320 0.000 1720.440 1.120 ;
 END
END DIA63
PIN DOA63
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1706.300 0.000 1707.420 1.120 ;
  LAYER metal4 ;
  RECT 1706.300 0.000 1707.420 1.120 ;
  LAYER metal3 ;
  RECT 1706.300 0.000 1707.420 1.120 ;
  LAYER metal2 ;
  RECT 1706.300 0.000 1707.420 1.120 ;
  LAYER metal1 ;
  RECT 1706.300 0.000 1707.420 1.120 ;
 END
END DOA63
PIN DIA62
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1692.660 0.000 1693.780 1.120 ;
  LAYER metal4 ;
  RECT 1692.660 0.000 1693.780 1.120 ;
  LAYER metal3 ;
  RECT 1692.660 0.000 1693.780 1.120 ;
  LAYER metal2 ;
  RECT 1692.660 0.000 1693.780 1.120 ;
  LAYER metal1 ;
  RECT 1692.660 0.000 1693.780 1.120 ;
 END
END DIA62
PIN DOA62
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1679.020 0.000 1680.140 1.120 ;
  LAYER metal4 ;
  RECT 1679.020 0.000 1680.140 1.120 ;
  LAYER metal3 ;
  RECT 1679.020 0.000 1680.140 1.120 ;
  LAYER metal2 ;
  RECT 1679.020 0.000 1680.140 1.120 ;
  LAYER metal1 ;
  RECT 1679.020 0.000 1680.140 1.120 ;
 END
END DOA62
PIN DIA61
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1666.000 0.000 1667.120 1.120 ;
  LAYER metal4 ;
  RECT 1666.000 0.000 1667.120 1.120 ;
  LAYER metal3 ;
  RECT 1666.000 0.000 1667.120 1.120 ;
  LAYER metal2 ;
  RECT 1666.000 0.000 1667.120 1.120 ;
  LAYER metal1 ;
  RECT 1666.000 0.000 1667.120 1.120 ;
 END
END DIA61
PIN DOA61
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1652.360 0.000 1653.480 1.120 ;
  LAYER metal4 ;
  RECT 1652.360 0.000 1653.480 1.120 ;
  LAYER metal3 ;
  RECT 1652.360 0.000 1653.480 1.120 ;
  LAYER metal2 ;
  RECT 1652.360 0.000 1653.480 1.120 ;
  LAYER metal1 ;
  RECT 1652.360 0.000 1653.480 1.120 ;
 END
END DOA61
PIN DIA60
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1638.720 0.000 1639.840 1.120 ;
  LAYER metal4 ;
  RECT 1638.720 0.000 1639.840 1.120 ;
  LAYER metal3 ;
  RECT 1638.720 0.000 1639.840 1.120 ;
  LAYER metal2 ;
  RECT 1638.720 0.000 1639.840 1.120 ;
  LAYER metal1 ;
  RECT 1638.720 0.000 1639.840 1.120 ;
 END
END DIA60
PIN DOA60
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1625.700 0.000 1626.820 1.120 ;
  LAYER metal4 ;
  RECT 1625.700 0.000 1626.820 1.120 ;
  LAYER metal3 ;
  RECT 1625.700 0.000 1626.820 1.120 ;
  LAYER metal2 ;
  RECT 1625.700 0.000 1626.820 1.120 ;
  LAYER metal1 ;
  RECT 1625.700 0.000 1626.820 1.120 ;
 END
END DOA60
PIN DIA59
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1612.060 0.000 1613.180 1.120 ;
  LAYER metal4 ;
  RECT 1612.060 0.000 1613.180 1.120 ;
  LAYER metal3 ;
  RECT 1612.060 0.000 1613.180 1.120 ;
  LAYER metal2 ;
  RECT 1612.060 0.000 1613.180 1.120 ;
  LAYER metal1 ;
  RECT 1612.060 0.000 1613.180 1.120 ;
 END
END DIA59
PIN DOA59
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1598.420 0.000 1599.540 1.120 ;
  LAYER metal4 ;
  RECT 1598.420 0.000 1599.540 1.120 ;
  LAYER metal3 ;
  RECT 1598.420 0.000 1599.540 1.120 ;
  LAYER metal2 ;
  RECT 1598.420 0.000 1599.540 1.120 ;
  LAYER metal1 ;
  RECT 1598.420 0.000 1599.540 1.120 ;
 END
END DOA59
PIN DIA58
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1585.400 0.000 1586.520 1.120 ;
  LAYER metal4 ;
  RECT 1585.400 0.000 1586.520 1.120 ;
  LAYER metal3 ;
  RECT 1585.400 0.000 1586.520 1.120 ;
  LAYER metal2 ;
  RECT 1585.400 0.000 1586.520 1.120 ;
  LAYER metal1 ;
  RECT 1585.400 0.000 1586.520 1.120 ;
 END
END DIA58
PIN DOA58
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1571.760 0.000 1572.880 1.120 ;
  LAYER metal4 ;
  RECT 1571.760 0.000 1572.880 1.120 ;
  LAYER metal3 ;
  RECT 1571.760 0.000 1572.880 1.120 ;
  LAYER metal2 ;
  RECT 1571.760 0.000 1572.880 1.120 ;
  LAYER metal1 ;
  RECT 1571.760 0.000 1572.880 1.120 ;
 END
END DOA58
PIN DIA57
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1558.120 0.000 1559.240 1.120 ;
  LAYER metal4 ;
  RECT 1558.120 0.000 1559.240 1.120 ;
  LAYER metal3 ;
  RECT 1558.120 0.000 1559.240 1.120 ;
  LAYER metal2 ;
  RECT 1558.120 0.000 1559.240 1.120 ;
  LAYER metal1 ;
  RECT 1558.120 0.000 1559.240 1.120 ;
 END
END DIA57
PIN DOA57
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1545.100 0.000 1546.220 1.120 ;
  LAYER metal4 ;
  RECT 1545.100 0.000 1546.220 1.120 ;
  LAYER metal3 ;
  RECT 1545.100 0.000 1546.220 1.120 ;
  LAYER metal2 ;
  RECT 1545.100 0.000 1546.220 1.120 ;
  LAYER metal1 ;
  RECT 1545.100 0.000 1546.220 1.120 ;
 END
END DOA57
PIN DIA56
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1531.460 0.000 1532.580 1.120 ;
  LAYER metal4 ;
  RECT 1531.460 0.000 1532.580 1.120 ;
  LAYER metal3 ;
  RECT 1531.460 0.000 1532.580 1.120 ;
  LAYER metal2 ;
  RECT 1531.460 0.000 1532.580 1.120 ;
  LAYER metal1 ;
  RECT 1531.460 0.000 1532.580 1.120 ;
 END
END DIA56
PIN DOA56
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1517.820 0.000 1518.940 1.120 ;
  LAYER metal4 ;
  RECT 1517.820 0.000 1518.940 1.120 ;
  LAYER metal3 ;
  RECT 1517.820 0.000 1518.940 1.120 ;
  LAYER metal2 ;
  RECT 1517.820 0.000 1518.940 1.120 ;
  LAYER metal1 ;
  RECT 1517.820 0.000 1518.940 1.120 ;
 END
END DOA56
PIN DIA55
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1504.800 0.000 1505.920 1.120 ;
  LAYER metal4 ;
  RECT 1504.800 0.000 1505.920 1.120 ;
  LAYER metal3 ;
  RECT 1504.800 0.000 1505.920 1.120 ;
  LAYER metal2 ;
  RECT 1504.800 0.000 1505.920 1.120 ;
  LAYER metal1 ;
  RECT 1504.800 0.000 1505.920 1.120 ;
 END
END DIA55
PIN DOA55
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1491.160 0.000 1492.280 1.120 ;
  LAYER metal4 ;
  RECT 1491.160 0.000 1492.280 1.120 ;
  LAYER metal3 ;
  RECT 1491.160 0.000 1492.280 1.120 ;
  LAYER metal2 ;
  RECT 1491.160 0.000 1492.280 1.120 ;
  LAYER metal1 ;
  RECT 1491.160 0.000 1492.280 1.120 ;
 END
END DOA55
PIN DIA54
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1477.520 0.000 1478.640 1.120 ;
  LAYER metal4 ;
  RECT 1477.520 0.000 1478.640 1.120 ;
  LAYER metal3 ;
  RECT 1477.520 0.000 1478.640 1.120 ;
  LAYER metal2 ;
  RECT 1477.520 0.000 1478.640 1.120 ;
  LAYER metal1 ;
  RECT 1477.520 0.000 1478.640 1.120 ;
 END
END DIA54
PIN DOA54
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1464.500 0.000 1465.620 1.120 ;
  LAYER metal4 ;
  RECT 1464.500 0.000 1465.620 1.120 ;
  LAYER metal3 ;
  RECT 1464.500 0.000 1465.620 1.120 ;
  LAYER metal2 ;
  RECT 1464.500 0.000 1465.620 1.120 ;
  LAYER metal1 ;
  RECT 1464.500 0.000 1465.620 1.120 ;
 END
END DOA54
PIN DIA53
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1450.860 0.000 1451.980 1.120 ;
  LAYER metal4 ;
  RECT 1450.860 0.000 1451.980 1.120 ;
  LAYER metal3 ;
  RECT 1450.860 0.000 1451.980 1.120 ;
  LAYER metal2 ;
  RECT 1450.860 0.000 1451.980 1.120 ;
  LAYER metal1 ;
  RECT 1450.860 0.000 1451.980 1.120 ;
 END
END DIA53
PIN DOA53
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1437.220 0.000 1438.340 1.120 ;
  LAYER metal4 ;
  RECT 1437.220 0.000 1438.340 1.120 ;
  LAYER metal3 ;
  RECT 1437.220 0.000 1438.340 1.120 ;
  LAYER metal2 ;
  RECT 1437.220 0.000 1438.340 1.120 ;
  LAYER metal1 ;
  RECT 1437.220 0.000 1438.340 1.120 ;
 END
END DOA53
PIN DIA52
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1424.200 0.000 1425.320 1.120 ;
  LAYER metal4 ;
  RECT 1424.200 0.000 1425.320 1.120 ;
  LAYER metal3 ;
  RECT 1424.200 0.000 1425.320 1.120 ;
  LAYER metal2 ;
  RECT 1424.200 0.000 1425.320 1.120 ;
  LAYER metal1 ;
  RECT 1424.200 0.000 1425.320 1.120 ;
 END
END DIA52
PIN DOA52
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1410.560 0.000 1411.680 1.120 ;
  LAYER metal4 ;
  RECT 1410.560 0.000 1411.680 1.120 ;
  LAYER metal3 ;
  RECT 1410.560 0.000 1411.680 1.120 ;
  LAYER metal2 ;
  RECT 1410.560 0.000 1411.680 1.120 ;
  LAYER metal1 ;
  RECT 1410.560 0.000 1411.680 1.120 ;
 END
END DOA52
PIN DIA51
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1396.920 0.000 1398.040 1.120 ;
  LAYER metal4 ;
  RECT 1396.920 0.000 1398.040 1.120 ;
  LAYER metal3 ;
  RECT 1396.920 0.000 1398.040 1.120 ;
  LAYER metal2 ;
  RECT 1396.920 0.000 1398.040 1.120 ;
  LAYER metal1 ;
  RECT 1396.920 0.000 1398.040 1.120 ;
 END
END DIA51
PIN DOA51
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1383.900 0.000 1385.020 1.120 ;
  LAYER metal4 ;
  RECT 1383.900 0.000 1385.020 1.120 ;
  LAYER metal3 ;
  RECT 1383.900 0.000 1385.020 1.120 ;
  LAYER metal2 ;
  RECT 1383.900 0.000 1385.020 1.120 ;
  LAYER metal1 ;
  RECT 1383.900 0.000 1385.020 1.120 ;
 END
END DOA51
PIN DIA50
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1370.260 0.000 1371.380 1.120 ;
  LAYER metal4 ;
  RECT 1370.260 0.000 1371.380 1.120 ;
  LAYER metal3 ;
  RECT 1370.260 0.000 1371.380 1.120 ;
  LAYER metal2 ;
  RECT 1370.260 0.000 1371.380 1.120 ;
  LAYER metal1 ;
  RECT 1370.260 0.000 1371.380 1.120 ;
 END
END DIA50
PIN DOA50
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1356.620 0.000 1357.740 1.120 ;
  LAYER metal4 ;
  RECT 1356.620 0.000 1357.740 1.120 ;
  LAYER metal3 ;
  RECT 1356.620 0.000 1357.740 1.120 ;
  LAYER metal2 ;
  RECT 1356.620 0.000 1357.740 1.120 ;
  LAYER metal1 ;
  RECT 1356.620 0.000 1357.740 1.120 ;
 END
END DOA50
PIN DIA49
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1343.600 0.000 1344.720 1.120 ;
  LAYER metal4 ;
  RECT 1343.600 0.000 1344.720 1.120 ;
  LAYER metal3 ;
  RECT 1343.600 0.000 1344.720 1.120 ;
  LAYER metal2 ;
  RECT 1343.600 0.000 1344.720 1.120 ;
  LAYER metal1 ;
  RECT 1343.600 0.000 1344.720 1.120 ;
 END
END DIA49
PIN DOA49
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1329.960 0.000 1331.080 1.120 ;
  LAYER metal4 ;
  RECT 1329.960 0.000 1331.080 1.120 ;
  LAYER metal3 ;
  RECT 1329.960 0.000 1331.080 1.120 ;
  LAYER metal2 ;
  RECT 1329.960 0.000 1331.080 1.120 ;
  LAYER metal1 ;
  RECT 1329.960 0.000 1331.080 1.120 ;
 END
END DOA49
PIN DIA48
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1316.320 0.000 1317.440 1.120 ;
  LAYER metal4 ;
  RECT 1316.320 0.000 1317.440 1.120 ;
  LAYER metal3 ;
  RECT 1316.320 0.000 1317.440 1.120 ;
  LAYER metal2 ;
  RECT 1316.320 0.000 1317.440 1.120 ;
  LAYER metal1 ;
  RECT 1316.320 0.000 1317.440 1.120 ;
 END
END DIA48
PIN DOA48
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1302.680 0.000 1303.800 1.120 ;
  LAYER metal4 ;
  RECT 1302.680 0.000 1303.800 1.120 ;
  LAYER metal3 ;
  RECT 1302.680 0.000 1303.800 1.120 ;
  LAYER metal2 ;
  RECT 1302.680 0.000 1303.800 1.120 ;
  LAYER metal1 ;
  RECT 1302.680 0.000 1303.800 1.120 ;
 END
END DOA48
PIN DIA47
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1289.660 0.000 1290.780 1.120 ;
  LAYER metal4 ;
  RECT 1289.660 0.000 1290.780 1.120 ;
  LAYER metal3 ;
  RECT 1289.660 0.000 1290.780 1.120 ;
  LAYER metal2 ;
  RECT 1289.660 0.000 1290.780 1.120 ;
  LAYER metal1 ;
  RECT 1289.660 0.000 1290.780 1.120 ;
 END
END DIA47
PIN DOA47
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1276.020 0.000 1277.140 1.120 ;
  LAYER metal4 ;
  RECT 1276.020 0.000 1277.140 1.120 ;
  LAYER metal3 ;
  RECT 1276.020 0.000 1277.140 1.120 ;
  LAYER metal2 ;
  RECT 1276.020 0.000 1277.140 1.120 ;
  LAYER metal1 ;
  RECT 1276.020 0.000 1277.140 1.120 ;
 END
END DOA47
PIN DIA46
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1262.380 0.000 1263.500 1.120 ;
  LAYER metal4 ;
  RECT 1262.380 0.000 1263.500 1.120 ;
  LAYER metal3 ;
  RECT 1262.380 0.000 1263.500 1.120 ;
  LAYER metal2 ;
  RECT 1262.380 0.000 1263.500 1.120 ;
  LAYER metal1 ;
  RECT 1262.380 0.000 1263.500 1.120 ;
 END
END DIA46
PIN DOA46
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1249.360 0.000 1250.480 1.120 ;
  LAYER metal4 ;
  RECT 1249.360 0.000 1250.480 1.120 ;
  LAYER metal3 ;
  RECT 1249.360 0.000 1250.480 1.120 ;
  LAYER metal2 ;
  RECT 1249.360 0.000 1250.480 1.120 ;
  LAYER metal1 ;
  RECT 1249.360 0.000 1250.480 1.120 ;
 END
END DOA46
PIN DIA45
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1235.720 0.000 1236.840 1.120 ;
  LAYER metal4 ;
  RECT 1235.720 0.000 1236.840 1.120 ;
  LAYER metal3 ;
  RECT 1235.720 0.000 1236.840 1.120 ;
  LAYER metal2 ;
  RECT 1235.720 0.000 1236.840 1.120 ;
  LAYER metal1 ;
  RECT 1235.720 0.000 1236.840 1.120 ;
 END
END DIA45
PIN DOA45
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1222.080 0.000 1223.200 1.120 ;
  LAYER metal4 ;
  RECT 1222.080 0.000 1223.200 1.120 ;
  LAYER metal3 ;
  RECT 1222.080 0.000 1223.200 1.120 ;
  LAYER metal2 ;
  RECT 1222.080 0.000 1223.200 1.120 ;
  LAYER metal1 ;
  RECT 1222.080 0.000 1223.200 1.120 ;
 END
END DOA45
PIN DIA44
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1209.060 0.000 1210.180 1.120 ;
  LAYER metal4 ;
  RECT 1209.060 0.000 1210.180 1.120 ;
  LAYER metal3 ;
  RECT 1209.060 0.000 1210.180 1.120 ;
  LAYER metal2 ;
  RECT 1209.060 0.000 1210.180 1.120 ;
  LAYER metal1 ;
  RECT 1209.060 0.000 1210.180 1.120 ;
 END
END DIA44
PIN DOA44
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1195.420 0.000 1196.540 1.120 ;
  LAYER metal4 ;
  RECT 1195.420 0.000 1196.540 1.120 ;
  LAYER metal3 ;
  RECT 1195.420 0.000 1196.540 1.120 ;
  LAYER metal2 ;
  RECT 1195.420 0.000 1196.540 1.120 ;
  LAYER metal1 ;
  RECT 1195.420 0.000 1196.540 1.120 ;
 END
END DOA44
PIN DIA43
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1181.780 0.000 1182.900 1.120 ;
  LAYER metal4 ;
  RECT 1181.780 0.000 1182.900 1.120 ;
  LAYER metal3 ;
  RECT 1181.780 0.000 1182.900 1.120 ;
  LAYER metal2 ;
  RECT 1181.780 0.000 1182.900 1.120 ;
  LAYER metal1 ;
  RECT 1181.780 0.000 1182.900 1.120 ;
 END
END DIA43
PIN DOA43
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1168.760 0.000 1169.880 1.120 ;
  LAYER metal4 ;
  RECT 1168.760 0.000 1169.880 1.120 ;
  LAYER metal3 ;
  RECT 1168.760 0.000 1169.880 1.120 ;
  LAYER metal2 ;
  RECT 1168.760 0.000 1169.880 1.120 ;
  LAYER metal1 ;
  RECT 1168.760 0.000 1169.880 1.120 ;
 END
END DOA43
PIN DIA42
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1155.120 0.000 1156.240 1.120 ;
  LAYER metal4 ;
  RECT 1155.120 0.000 1156.240 1.120 ;
  LAYER metal3 ;
  RECT 1155.120 0.000 1156.240 1.120 ;
  LAYER metal2 ;
  RECT 1155.120 0.000 1156.240 1.120 ;
  LAYER metal1 ;
  RECT 1155.120 0.000 1156.240 1.120 ;
 END
END DIA42
PIN DOA42
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1141.480 0.000 1142.600 1.120 ;
  LAYER metal4 ;
  RECT 1141.480 0.000 1142.600 1.120 ;
  LAYER metal3 ;
  RECT 1141.480 0.000 1142.600 1.120 ;
  LAYER metal2 ;
  RECT 1141.480 0.000 1142.600 1.120 ;
  LAYER metal1 ;
  RECT 1141.480 0.000 1142.600 1.120 ;
 END
END DOA42
PIN DIA41
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1128.460 0.000 1129.580 1.120 ;
  LAYER metal4 ;
  RECT 1128.460 0.000 1129.580 1.120 ;
  LAYER metal3 ;
  RECT 1128.460 0.000 1129.580 1.120 ;
  LAYER metal2 ;
  RECT 1128.460 0.000 1129.580 1.120 ;
  LAYER metal1 ;
  RECT 1128.460 0.000 1129.580 1.120 ;
 END
END DIA41
PIN DOA41
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1114.820 0.000 1115.940 1.120 ;
  LAYER metal4 ;
  RECT 1114.820 0.000 1115.940 1.120 ;
  LAYER metal3 ;
  RECT 1114.820 0.000 1115.940 1.120 ;
  LAYER metal2 ;
  RECT 1114.820 0.000 1115.940 1.120 ;
  LAYER metal1 ;
  RECT 1114.820 0.000 1115.940 1.120 ;
 END
END DOA41
PIN DIA40
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1101.180 0.000 1102.300 1.120 ;
  LAYER metal4 ;
  RECT 1101.180 0.000 1102.300 1.120 ;
  LAYER metal3 ;
  RECT 1101.180 0.000 1102.300 1.120 ;
  LAYER metal2 ;
  RECT 1101.180 0.000 1102.300 1.120 ;
  LAYER metal1 ;
  RECT 1101.180 0.000 1102.300 1.120 ;
 END
END DIA40
PIN DOA40
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1088.160 0.000 1089.280 1.120 ;
  LAYER metal4 ;
  RECT 1088.160 0.000 1089.280 1.120 ;
  LAYER metal3 ;
  RECT 1088.160 0.000 1089.280 1.120 ;
  LAYER metal2 ;
  RECT 1088.160 0.000 1089.280 1.120 ;
  LAYER metal1 ;
  RECT 1088.160 0.000 1089.280 1.120 ;
 END
END DOA40
PIN DIA39
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 1074.520 0.000 1075.640 1.120 ;
  LAYER metal4 ;
  RECT 1074.520 0.000 1075.640 1.120 ;
  LAYER metal3 ;
  RECT 1074.520 0.000 1075.640 1.120 ;
  LAYER metal2 ;
  RECT 1074.520 0.000 1075.640 1.120 ;
  LAYER metal1 ;
  RECT 1074.520 0.000 1075.640 1.120 ;
 END
END DIA39
PIN DOA39
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1060.880 0.000 1062.000 1.120 ;
  LAYER metal4 ;
  RECT 1060.880 0.000 1062.000 1.120 ;
  LAYER metal3 ;
  RECT 1060.880 0.000 1062.000 1.120 ;
  LAYER metal2 ;
  RECT 1060.880 0.000 1062.000 1.120 ;
  LAYER metal1 ;
  RECT 1060.880 0.000 1062.000 1.120 ;
 END
END DOA39
PIN DIA38
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1047.860 0.000 1048.980 1.120 ;
  LAYER metal4 ;
  RECT 1047.860 0.000 1048.980 1.120 ;
  LAYER metal3 ;
  RECT 1047.860 0.000 1048.980 1.120 ;
  LAYER metal2 ;
  RECT 1047.860 0.000 1048.980 1.120 ;
  LAYER metal1 ;
  RECT 1047.860 0.000 1048.980 1.120 ;
 END
END DIA38
PIN DOA38
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 1034.220 0.000 1035.340 1.120 ;
  LAYER metal4 ;
  RECT 1034.220 0.000 1035.340 1.120 ;
  LAYER metal3 ;
  RECT 1034.220 0.000 1035.340 1.120 ;
  LAYER metal2 ;
  RECT 1034.220 0.000 1035.340 1.120 ;
  LAYER metal1 ;
  RECT 1034.220 0.000 1035.340 1.120 ;
 END
END DOA38
PIN DIA37
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 1020.580 0.000 1021.700 1.120 ;
  LAYER metal4 ;
  RECT 1020.580 0.000 1021.700 1.120 ;
  LAYER metal3 ;
  RECT 1020.580 0.000 1021.700 1.120 ;
  LAYER metal2 ;
  RECT 1020.580 0.000 1021.700 1.120 ;
  LAYER metal1 ;
  RECT 1020.580 0.000 1021.700 1.120 ;
 END
END DIA37
PIN DOA37
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 1007.560 0.000 1008.680 1.120 ;
  LAYER metal4 ;
  RECT 1007.560 0.000 1008.680 1.120 ;
  LAYER metal3 ;
  RECT 1007.560 0.000 1008.680 1.120 ;
  LAYER metal2 ;
  RECT 1007.560 0.000 1008.680 1.120 ;
  LAYER metal1 ;
  RECT 1007.560 0.000 1008.680 1.120 ;
 END
END DOA37
PIN DIA36
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 993.920 0.000 995.040 1.120 ;
  LAYER metal4 ;
  RECT 993.920 0.000 995.040 1.120 ;
  LAYER metal3 ;
  RECT 993.920 0.000 995.040 1.120 ;
  LAYER metal2 ;
  RECT 993.920 0.000 995.040 1.120 ;
  LAYER metal1 ;
  RECT 993.920 0.000 995.040 1.120 ;
 END
END DIA36
PIN DOA36
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 980.280 0.000 981.400 1.120 ;
  LAYER metal4 ;
  RECT 980.280 0.000 981.400 1.120 ;
  LAYER metal3 ;
  RECT 980.280 0.000 981.400 1.120 ;
  LAYER metal2 ;
  RECT 980.280 0.000 981.400 1.120 ;
  LAYER metal1 ;
  RECT 980.280 0.000 981.400 1.120 ;
 END
END DOA36
PIN DIA35
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 967.260 0.000 968.380 1.120 ;
  LAYER metal4 ;
  RECT 967.260 0.000 968.380 1.120 ;
  LAYER metal3 ;
  RECT 967.260 0.000 968.380 1.120 ;
  LAYER metal2 ;
  RECT 967.260 0.000 968.380 1.120 ;
  LAYER metal1 ;
  RECT 967.260 0.000 968.380 1.120 ;
 END
END DIA35
PIN DOA35
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 953.620 0.000 954.740 1.120 ;
  LAYER metal4 ;
  RECT 953.620 0.000 954.740 1.120 ;
  LAYER metal3 ;
  RECT 953.620 0.000 954.740 1.120 ;
  LAYER metal2 ;
  RECT 953.620 0.000 954.740 1.120 ;
  LAYER metal1 ;
  RECT 953.620 0.000 954.740 1.120 ;
 END
END DOA35
PIN DIA34
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 939.980 0.000 941.100 1.120 ;
  LAYER metal4 ;
  RECT 939.980 0.000 941.100 1.120 ;
  LAYER metal3 ;
  RECT 939.980 0.000 941.100 1.120 ;
  LAYER metal2 ;
  RECT 939.980 0.000 941.100 1.120 ;
  LAYER metal1 ;
  RECT 939.980 0.000 941.100 1.120 ;
 END
END DIA34
PIN DOA34
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 926.960 0.000 928.080 1.120 ;
  LAYER metal4 ;
  RECT 926.960 0.000 928.080 1.120 ;
  LAYER metal3 ;
  RECT 926.960 0.000 928.080 1.120 ;
  LAYER metal2 ;
  RECT 926.960 0.000 928.080 1.120 ;
  LAYER metal1 ;
  RECT 926.960 0.000 928.080 1.120 ;
 END
END DOA34
PIN DIA33
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 913.320 0.000 914.440 1.120 ;
  LAYER metal4 ;
  RECT 913.320 0.000 914.440 1.120 ;
  LAYER metal3 ;
  RECT 913.320 0.000 914.440 1.120 ;
  LAYER metal2 ;
  RECT 913.320 0.000 914.440 1.120 ;
  LAYER metal1 ;
  RECT 913.320 0.000 914.440 1.120 ;
 END
END DIA33
PIN DOA33
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 899.680 0.000 900.800 1.120 ;
  LAYER metal4 ;
  RECT 899.680 0.000 900.800 1.120 ;
  LAYER metal3 ;
  RECT 899.680 0.000 900.800 1.120 ;
  LAYER metal2 ;
  RECT 899.680 0.000 900.800 1.120 ;
  LAYER metal1 ;
  RECT 899.680 0.000 900.800 1.120 ;
 END
END DOA33
PIN DIA32
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 886.040 0.000 887.160 1.120 ;
  LAYER metal4 ;
  RECT 886.040 0.000 887.160 1.120 ;
  LAYER metal3 ;
  RECT 886.040 0.000 887.160 1.120 ;
  LAYER metal2 ;
  RECT 886.040 0.000 887.160 1.120 ;
  LAYER metal1 ;
  RECT 886.040 0.000 887.160 1.120 ;
 END
END DIA32
PIN DOA32
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 873.020 0.000 874.140 1.120 ;
  LAYER metal4 ;
  RECT 873.020 0.000 874.140 1.120 ;
  LAYER metal3 ;
  RECT 873.020 0.000 874.140 1.120 ;
  LAYER metal2 ;
  RECT 873.020 0.000 874.140 1.120 ;
  LAYER metal1 ;
  RECT 873.020 0.000 874.140 1.120 ;
 END
END DOA32
PIN DIA31
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 859.380 0.000 860.500 1.120 ;
  LAYER metal4 ;
  RECT 859.380 0.000 860.500 1.120 ;
  LAYER metal3 ;
  RECT 859.380 0.000 860.500 1.120 ;
  LAYER metal2 ;
  RECT 859.380 0.000 860.500 1.120 ;
  LAYER metal1 ;
  RECT 859.380 0.000 860.500 1.120 ;
 END
END DIA31
PIN DOA31
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 845.740 0.000 846.860 1.120 ;
  LAYER metal4 ;
  RECT 845.740 0.000 846.860 1.120 ;
  LAYER metal3 ;
  RECT 845.740 0.000 846.860 1.120 ;
  LAYER metal2 ;
  RECT 845.740 0.000 846.860 1.120 ;
  LAYER metal1 ;
  RECT 845.740 0.000 846.860 1.120 ;
 END
END DOA31
PIN DIA30
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 832.720 0.000 833.840 1.120 ;
  LAYER metal4 ;
  RECT 832.720 0.000 833.840 1.120 ;
  LAYER metal3 ;
  RECT 832.720 0.000 833.840 1.120 ;
  LAYER metal2 ;
  RECT 832.720 0.000 833.840 1.120 ;
  LAYER metal1 ;
  RECT 832.720 0.000 833.840 1.120 ;
 END
END DIA30
PIN DOA30
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 819.080 0.000 820.200 1.120 ;
  LAYER metal4 ;
  RECT 819.080 0.000 820.200 1.120 ;
  LAYER metal3 ;
  RECT 819.080 0.000 820.200 1.120 ;
  LAYER metal2 ;
  RECT 819.080 0.000 820.200 1.120 ;
  LAYER metal1 ;
  RECT 819.080 0.000 820.200 1.120 ;
 END
END DOA30
PIN DIA29
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 805.440 0.000 806.560 1.120 ;
  LAYER metal4 ;
  RECT 805.440 0.000 806.560 1.120 ;
  LAYER metal3 ;
  RECT 805.440 0.000 806.560 1.120 ;
  LAYER metal2 ;
  RECT 805.440 0.000 806.560 1.120 ;
  LAYER metal1 ;
  RECT 805.440 0.000 806.560 1.120 ;
 END
END DIA29
PIN DOA29
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 792.420 0.000 793.540 1.120 ;
  LAYER metal4 ;
  RECT 792.420 0.000 793.540 1.120 ;
  LAYER metal3 ;
  RECT 792.420 0.000 793.540 1.120 ;
  LAYER metal2 ;
  RECT 792.420 0.000 793.540 1.120 ;
  LAYER metal1 ;
  RECT 792.420 0.000 793.540 1.120 ;
 END
END DOA29
PIN DIA28
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 778.780 0.000 779.900 1.120 ;
  LAYER metal4 ;
  RECT 778.780 0.000 779.900 1.120 ;
  LAYER metal3 ;
  RECT 778.780 0.000 779.900 1.120 ;
  LAYER metal2 ;
  RECT 778.780 0.000 779.900 1.120 ;
  LAYER metal1 ;
  RECT 778.780 0.000 779.900 1.120 ;
 END
END DIA28
PIN DOA28
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 765.140 0.000 766.260 1.120 ;
  LAYER metal4 ;
  RECT 765.140 0.000 766.260 1.120 ;
  LAYER metal3 ;
  RECT 765.140 0.000 766.260 1.120 ;
  LAYER metal2 ;
  RECT 765.140 0.000 766.260 1.120 ;
  LAYER metal1 ;
  RECT 765.140 0.000 766.260 1.120 ;
 END
END DOA28
PIN DIA27
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 752.120 0.000 753.240 1.120 ;
  LAYER metal4 ;
  RECT 752.120 0.000 753.240 1.120 ;
  LAYER metal3 ;
  RECT 752.120 0.000 753.240 1.120 ;
  LAYER metal2 ;
  RECT 752.120 0.000 753.240 1.120 ;
  LAYER metal1 ;
  RECT 752.120 0.000 753.240 1.120 ;
 END
END DIA27
PIN DOA27
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 738.480 0.000 739.600 1.120 ;
  LAYER metal4 ;
  RECT 738.480 0.000 739.600 1.120 ;
  LAYER metal3 ;
  RECT 738.480 0.000 739.600 1.120 ;
  LAYER metal2 ;
  RECT 738.480 0.000 739.600 1.120 ;
  LAYER metal1 ;
  RECT 738.480 0.000 739.600 1.120 ;
 END
END DOA27
PIN DIA26
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 724.840 0.000 725.960 1.120 ;
  LAYER metal4 ;
  RECT 724.840 0.000 725.960 1.120 ;
  LAYER metal3 ;
  RECT 724.840 0.000 725.960 1.120 ;
  LAYER metal2 ;
  RECT 724.840 0.000 725.960 1.120 ;
  LAYER metal1 ;
  RECT 724.840 0.000 725.960 1.120 ;
 END
END DIA26
PIN DOA26
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 711.820 0.000 712.940 1.120 ;
  LAYER metal4 ;
  RECT 711.820 0.000 712.940 1.120 ;
  LAYER metal3 ;
  RECT 711.820 0.000 712.940 1.120 ;
  LAYER metal2 ;
  RECT 711.820 0.000 712.940 1.120 ;
  LAYER metal1 ;
  RECT 711.820 0.000 712.940 1.120 ;
 END
END DOA26
PIN DIA25
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 698.180 0.000 699.300 1.120 ;
  LAYER metal4 ;
  RECT 698.180 0.000 699.300 1.120 ;
  LAYER metal3 ;
  RECT 698.180 0.000 699.300 1.120 ;
  LAYER metal2 ;
  RECT 698.180 0.000 699.300 1.120 ;
  LAYER metal1 ;
  RECT 698.180 0.000 699.300 1.120 ;
 END
END DIA25
PIN DOA25
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 684.540 0.000 685.660 1.120 ;
  LAYER metal4 ;
  RECT 684.540 0.000 685.660 1.120 ;
  LAYER metal3 ;
  RECT 684.540 0.000 685.660 1.120 ;
  LAYER metal2 ;
  RECT 684.540 0.000 685.660 1.120 ;
  LAYER metal1 ;
  RECT 684.540 0.000 685.660 1.120 ;
 END
END DOA25
PIN DIA24
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 671.520 0.000 672.640 1.120 ;
  LAYER metal4 ;
  RECT 671.520 0.000 672.640 1.120 ;
  LAYER metal3 ;
  RECT 671.520 0.000 672.640 1.120 ;
  LAYER metal2 ;
  RECT 671.520 0.000 672.640 1.120 ;
  LAYER metal1 ;
  RECT 671.520 0.000 672.640 1.120 ;
 END
END DIA24
PIN DOA24
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 657.880 0.000 659.000 1.120 ;
  LAYER metal4 ;
  RECT 657.880 0.000 659.000 1.120 ;
  LAYER metal3 ;
  RECT 657.880 0.000 659.000 1.120 ;
  LAYER metal2 ;
  RECT 657.880 0.000 659.000 1.120 ;
  LAYER metal1 ;
  RECT 657.880 0.000 659.000 1.120 ;
 END
END DOA24
PIN DIA23
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 644.240 0.000 645.360 1.120 ;
  LAYER metal4 ;
  RECT 644.240 0.000 645.360 1.120 ;
  LAYER metal3 ;
  RECT 644.240 0.000 645.360 1.120 ;
  LAYER metal2 ;
  RECT 644.240 0.000 645.360 1.120 ;
  LAYER metal1 ;
  RECT 644.240 0.000 645.360 1.120 ;
 END
END DIA23
PIN DOA23
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 631.220 0.000 632.340 1.120 ;
  LAYER metal4 ;
  RECT 631.220 0.000 632.340 1.120 ;
  LAYER metal3 ;
  RECT 631.220 0.000 632.340 1.120 ;
  LAYER metal2 ;
  RECT 631.220 0.000 632.340 1.120 ;
  LAYER metal1 ;
  RECT 631.220 0.000 632.340 1.120 ;
 END
END DOA23
PIN DIA22
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 617.580 0.000 618.700 1.120 ;
  LAYER metal4 ;
  RECT 617.580 0.000 618.700 1.120 ;
  LAYER metal3 ;
  RECT 617.580 0.000 618.700 1.120 ;
  LAYER metal2 ;
  RECT 617.580 0.000 618.700 1.120 ;
  LAYER metal1 ;
  RECT 617.580 0.000 618.700 1.120 ;
 END
END DIA22
PIN DOA22
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 603.940 0.000 605.060 1.120 ;
  LAYER metal4 ;
  RECT 603.940 0.000 605.060 1.120 ;
  LAYER metal3 ;
  RECT 603.940 0.000 605.060 1.120 ;
  LAYER metal2 ;
  RECT 603.940 0.000 605.060 1.120 ;
  LAYER metal1 ;
  RECT 603.940 0.000 605.060 1.120 ;
 END
END DOA22
PIN DIA21
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 590.920 0.000 592.040 1.120 ;
  LAYER metal4 ;
  RECT 590.920 0.000 592.040 1.120 ;
  LAYER metal3 ;
  RECT 590.920 0.000 592.040 1.120 ;
  LAYER metal2 ;
  RECT 590.920 0.000 592.040 1.120 ;
  LAYER metal1 ;
  RECT 590.920 0.000 592.040 1.120 ;
 END
END DIA21
PIN DOA21
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 577.280 0.000 578.400 1.120 ;
  LAYER metal4 ;
  RECT 577.280 0.000 578.400 1.120 ;
  LAYER metal3 ;
  RECT 577.280 0.000 578.400 1.120 ;
  LAYER metal2 ;
  RECT 577.280 0.000 578.400 1.120 ;
  LAYER metal1 ;
  RECT 577.280 0.000 578.400 1.120 ;
 END
END DOA21
PIN DIA20
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 563.640 0.000 564.760 1.120 ;
  LAYER metal4 ;
  RECT 563.640 0.000 564.760 1.120 ;
  LAYER metal3 ;
  RECT 563.640 0.000 564.760 1.120 ;
  LAYER metal2 ;
  RECT 563.640 0.000 564.760 1.120 ;
  LAYER metal1 ;
  RECT 563.640 0.000 564.760 1.120 ;
 END
END DIA20
PIN DOA20
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 550.620 0.000 551.740 1.120 ;
  LAYER metal4 ;
  RECT 550.620 0.000 551.740 1.120 ;
  LAYER metal3 ;
  RECT 550.620 0.000 551.740 1.120 ;
  LAYER metal2 ;
  RECT 550.620 0.000 551.740 1.120 ;
  LAYER metal1 ;
  RECT 550.620 0.000 551.740 1.120 ;
 END
END DOA20
PIN DIA19
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 536.980 0.000 538.100 1.120 ;
  LAYER metal4 ;
  RECT 536.980 0.000 538.100 1.120 ;
  LAYER metal3 ;
  RECT 536.980 0.000 538.100 1.120 ;
  LAYER metal2 ;
  RECT 536.980 0.000 538.100 1.120 ;
  LAYER metal1 ;
  RECT 536.980 0.000 538.100 1.120 ;
 END
END DIA19
PIN DOA19
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 523.340 0.000 524.460 1.120 ;
  LAYER metal4 ;
  RECT 523.340 0.000 524.460 1.120 ;
  LAYER metal3 ;
  RECT 523.340 0.000 524.460 1.120 ;
  LAYER metal2 ;
  RECT 523.340 0.000 524.460 1.120 ;
  LAYER metal1 ;
  RECT 523.340 0.000 524.460 1.120 ;
 END
END DOA19
PIN DIA18
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 510.320 0.000 511.440 1.120 ;
  LAYER metal4 ;
  RECT 510.320 0.000 511.440 1.120 ;
  LAYER metal3 ;
  RECT 510.320 0.000 511.440 1.120 ;
  LAYER metal2 ;
  RECT 510.320 0.000 511.440 1.120 ;
  LAYER metal1 ;
  RECT 510.320 0.000 511.440 1.120 ;
 END
END DIA18
PIN DOA18
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 496.680 0.000 497.800 1.120 ;
  LAYER metal4 ;
  RECT 496.680 0.000 497.800 1.120 ;
  LAYER metal3 ;
  RECT 496.680 0.000 497.800 1.120 ;
  LAYER metal2 ;
  RECT 496.680 0.000 497.800 1.120 ;
  LAYER metal1 ;
  RECT 496.680 0.000 497.800 1.120 ;
 END
END DOA18
PIN DIA17
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 483.040 0.000 484.160 1.120 ;
  LAYER metal4 ;
  RECT 483.040 0.000 484.160 1.120 ;
  LAYER metal3 ;
  RECT 483.040 0.000 484.160 1.120 ;
  LAYER metal2 ;
  RECT 483.040 0.000 484.160 1.120 ;
  LAYER metal1 ;
  RECT 483.040 0.000 484.160 1.120 ;
 END
END DIA17
PIN DOA17
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 469.400 0.000 470.520 1.120 ;
  LAYER metal4 ;
  RECT 469.400 0.000 470.520 1.120 ;
  LAYER metal3 ;
  RECT 469.400 0.000 470.520 1.120 ;
  LAYER metal2 ;
  RECT 469.400 0.000 470.520 1.120 ;
  LAYER metal1 ;
  RECT 469.400 0.000 470.520 1.120 ;
 END
END DOA17
PIN DIA16
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 456.380 0.000 457.500 1.120 ;
  LAYER metal4 ;
  RECT 456.380 0.000 457.500 1.120 ;
  LAYER metal3 ;
  RECT 456.380 0.000 457.500 1.120 ;
  LAYER metal2 ;
  RECT 456.380 0.000 457.500 1.120 ;
  LAYER metal1 ;
  RECT 456.380 0.000 457.500 1.120 ;
 END
END DIA16
PIN DOA16
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 442.740 0.000 443.860 1.120 ;
  LAYER metal4 ;
  RECT 442.740 0.000 443.860 1.120 ;
  LAYER metal3 ;
  RECT 442.740 0.000 443.860 1.120 ;
  LAYER metal2 ;
  RECT 442.740 0.000 443.860 1.120 ;
  LAYER metal1 ;
  RECT 442.740 0.000 443.860 1.120 ;
 END
END DOA16
PIN DIA15
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER metal4 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER metal3 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER metal2 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER metal1 ;
  RECT 429.100 0.000 430.220 1.120 ;
 END
END DIA15
PIN DOA15
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 416.080 0.000 417.200 1.120 ;
  LAYER metal4 ;
  RECT 416.080 0.000 417.200 1.120 ;
  LAYER metal3 ;
  RECT 416.080 0.000 417.200 1.120 ;
  LAYER metal2 ;
  RECT 416.080 0.000 417.200 1.120 ;
  LAYER metal1 ;
  RECT 416.080 0.000 417.200 1.120 ;
 END
END DOA15
PIN DIA14
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER metal4 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER metal3 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER metal2 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER metal1 ;
  RECT 402.440 0.000 403.560 1.120 ;
 END
END DIA14
PIN DOA14
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 388.800 0.000 389.920 1.120 ;
  LAYER metal4 ;
  RECT 388.800 0.000 389.920 1.120 ;
  LAYER metal3 ;
  RECT 388.800 0.000 389.920 1.120 ;
  LAYER metal2 ;
  RECT 388.800 0.000 389.920 1.120 ;
  LAYER metal1 ;
  RECT 388.800 0.000 389.920 1.120 ;
 END
END DOA14
PIN DIA13
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 375.780 0.000 376.900 1.120 ;
  LAYER metal4 ;
  RECT 375.780 0.000 376.900 1.120 ;
  LAYER metal3 ;
  RECT 375.780 0.000 376.900 1.120 ;
  LAYER metal2 ;
  RECT 375.780 0.000 376.900 1.120 ;
  LAYER metal1 ;
  RECT 375.780 0.000 376.900 1.120 ;
 END
END DIA13
PIN DOA13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 362.140 0.000 363.260 1.120 ;
  LAYER metal4 ;
  RECT 362.140 0.000 363.260 1.120 ;
  LAYER metal3 ;
  RECT 362.140 0.000 363.260 1.120 ;
  LAYER metal2 ;
  RECT 362.140 0.000 363.260 1.120 ;
  LAYER metal1 ;
  RECT 362.140 0.000 363.260 1.120 ;
 END
END DOA13
PIN DIA12
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 348.500 0.000 349.620 1.120 ;
  LAYER metal4 ;
  RECT 348.500 0.000 349.620 1.120 ;
  LAYER metal3 ;
  RECT 348.500 0.000 349.620 1.120 ;
  LAYER metal2 ;
  RECT 348.500 0.000 349.620 1.120 ;
  LAYER metal1 ;
  RECT 348.500 0.000 349.620 1.120 ;
 END
END DIA12
PIN DOA12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 335.480 0.000 336.600 1.120 ;
  LAYER metal4 ;
  RECT 335.480 0.000 336.600 1.120 ;
  LAYER metal3 ;
  RECT 335.480 0.000 336.600 1.120 ;
  LAYER metal2 ;
  RECT 335.480 0.000 336.600 1.120 ;
  LAYER metal1 ;
  RECT 335.480 0.000 336.600 1.120 ;
 END
END DOA12
PIN DIA11
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 321.840 0.000 322.960 1.120 ;
  LAYER metal4 ;
  RECT 321.840 0.000 322.960 1.120 ;
  LAYER metal3 ;
  RECT 321.840 0.000 322.960 1.120 ;
  LAYER metal2 ;
  RECT 321.840 0.000 322.960 1.120 ;
  LAYER metal1 ;
  RECT 321.840 0.000 322.960 1.120 ;
 END
END DIA11
PIN DOA11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 308.200 0.000 309.320 1.120 ;
  LAYER metal4 ;
  RECT 308.200 0.000 309.320 1.120 ;
  LAYER metal3 ;
  RECT 308.200 0.000 309.320 1.120 ;
  LAYER metal2 ;
  RECT 308.200 0.000 309.320 1.120 ;
  LAYER metal1 ;
  RECT 308.200 0.000 309.320 1.120 ;
 END
END DOA11
PIN DIA10
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 295.180 0.000 296.300 1.120 ;
  LAYER metal4 ;
  RECT 295.180 0.000 296.300 1.120 ;
  LAYER metal3 ;
  RECT 295.180 0.000 296.300 1.120 ;
  LAYER metal2 ;
  RECT 295.180 0.000 296.300 1.120 ;
  LAYER metal1 ;
  RECT 295.180 0.000 296.300 1.120 ;
 END
END DIA10
PIN DOA10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 281.540 0.000 282.660 1.120 ;
  LAYER metal4 ;
  RECT 281.540 0.000 282.660 1.120 ;
  LAYER metal3 ;
  RECT 281.540 0.000 282.660 1.120 ;
  LAYER metal2 ;
  RECT 281.540 0.000 282.660 1.120 ;
  LAYER metal1 ;
  RECT 281.540 0.000 282.660 1.120 ;
 END
END DOA10
PIN DIA9
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER metal4 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER metal3 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER metal2 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER metal1 ;
  RECT 267.900 0.000 269.020 1.120 ;
 END
END DIA9
PIN DOA9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER metal4 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER metal3 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER metal2 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER metal1 ;
  RECT 254.880 0.000 256.000 1.120 ;
 END
END DOA9
PIN DIA8
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER metal4 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER metal3 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER metal2 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER metal1 ;
  RECT 241.240 0.000 242.360 1.120 ;
 END
END DIA8
PIN DOA8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 227.600 0.000 228.720 1.120 ;
  LAYER metal4 ;
  RECT 227.600 0.000 228.720 1.120 ;
  LAYER metal3 ;
  RECT 227.600 0.000 228.720 1.120 ;
  LAYER metal2 ;
  RECT 227.600 0.000 228.720 1.120 ;
  LAYER metal1 ;
  RECT 227.600 0.000 228.720 1.120 ;
 END
END DOA8
PIN DIA7
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 214.580 0.000 215.700 1.120 ;
  LAYER metal4 ;
  RECT 214.580 0.000 215.700 1.120 ;
  LAYER metal3 ;
  RECT 214.580 0.000 215.700 1.120 ;
  LAYER metal2 ;
  RECT 214.580 0.000 215.700 1.120 ;
  LAYER metal1 ;
  RECT 214.580 0.000 215.700 1.120 ;
 END
END DIA7
PIN DOA7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 200.940 0.000 202.060 1.120 ;
  LAYER metal4 ;
  RECT 200.940 0.000 202.060 1.120 ;
  LAYER metal3 ;
  RECT 200.940 0.000 202.060 1.120 ;
  LAYER metal2 ;
  RECT 200.940 0.000 202.060 1.120 ;
  LAYER metal1 ;
  RECT 200.940 0.000 202.060 1.120 ;
 END
END DOA7
PIN DIA6
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER metal4 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER metal3 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER metal2 ;
  RECT 187.300 0.000 188.420 1.120 ;
  LAYER metal1 ;
  RECT 187.300 0.000 188.420 1.120 ;
 END
END DIA6
PIN DOA6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 174.280 0.000 175.400 1.120 ;
  LAYER metal4 ;
  RECT 174.280 0.000 175.400 1.120 ;
  LAYER metal3 ;
  RECT 174.280 0.000 175.400 1.120 ;
  LAYER metal2 ;
  RECT 174.280 0.000 175.400 1.120 ;
  LAYER metal1 ;
  RECT 174.280 0.000 175.400 1.120 ;
 END
END DOA6
PIN DIA5
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 160.640 0.000 161.760 1.120 ;
  LAYER metal4 ;
  RECT 160.640 0.000 161.760 1.120 ;
  LAYER metal3 ;
  RECT 160.640 0.000 161.760 1.120 ;
  LAYER metal2 ;
  RECT 160.640 0.000 161.760 1.120 ;
  LAYER metal1 ;
  RECT 160.640 0.000 161.760 1.120 ;
 END
END DIA5
PIN DOA5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 147.000 0.000 148.120 1.120 ;
  LAYER metal4 ;
  RECT 147.000 0.000 148.120 1.120 ;
  LAYER metal3 ;
  RECT 147.000 0.000 148.120 1.120 ;
  LAYER metal2 ;
  RECT 147.000 0.000 148.120 1.120 ;
  LAYER metal1 ;
  RECT 147.000 0.000 148.120 1.120 ;
 END
END DOA5
PIN DIA4
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 133.980 0.000 135.100 1.120 ;
  LAYER metal4 ;
  RECT 133.980 0.000 135.100 1.120 ;
  LAYER metal3 ;
  RECT 133.980 0.000 135.100 1.120 ;
  LAYER metal2 ;
  RECT 133.980 0.000 135.100 1.120 ;
  LAYER metal1 ;
  RECT 133.980 0.000 135.100 1.120 ;
 END
END DIA4
PIN DOA4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 120.340 0.000 121.460 1.120 ;
  LAYER metal4 ;
  RECT 120.340 0.000 121.460 1.120 ;
  LAYER metal3 ;
  RECT 120.340 0.000 121.460 1.120 ;
  LAYER metal2 ;
  RECT 120.340 0.000 121.460 1.120 ;
  LAYER metal1 ;
  RECT 120.340 0.000 121.460 1.120 ;
 END
END DOA4
PIN DIA3
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal4 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal3 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal2 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal1 ;
  RECT 106.700 0.000 107.820 1.120 ;
 END
END DIA3
PIN DOA3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 93.680 0.000 94.800 1.120 ;
  LAYER metal4 ;
  RECT 93.680 0.000 94.800 1.120 ;
  LAYER metal3 ;
  RECT 93.680 0.000 94.800 1.120 ;
  LAYER metal2 ;
  RECT 93.680 0.000 94.800 1.120 ;
  LAYER metal1 ;
  RECT 93.680 0.000 94.800 1.120 ;
 END
END DOA3
PIN DIA2
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 80.040 0.000 81.160 1.120 ;
  LAYER metal4 ;
  RECT 80.040 0.000 81.160 1.120 ;
  LAYER metal3 ;
  RECT 80.040 0.000 81.160 1.120 ;
  LAYER metal2 ;
  RECT 80.040 0.000 81.160 1.120 ;
  LAYER metal1 ;
  RECT 80.040 0.000 81.160 1.120 ;
 END
END DIA2
PIN DOA2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 66.400 0.000 67.520 1.120 ;
  LAYER metal4 ;
  RECT 66.400 0.000 67.520 1.120 ;
  LAYER metal3 ;
  RECT 66.400 0.000 67.520 1.120 ;
  LAYER metal2 ;
  RECT 66.400 0.000 67.520 1.120 ;
  LAYER metal1 ;
  RECT 66.400 0.000 67.520 1.120 ;
 END
END DOA2
PIN DIA1
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal5 ;
  RECT 52.760 0.000 53.880 1.120 ;
  LAYER metal4 ;
  RECT 52.760 0.000 53.880 1.120 ;
  LAYER metal3 ;
  RECT 52.760 0.000 53.880 1.120 ;
  LAYER metal2 ;
  RECT 52.760 0.000 53.880 1.120 ;
  LAYER metal1 ;
  RECT 52.760 0.000 53.880 1.120 ;
 END
END DIA1
PIN DOA1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal5 ;
  RECT 39.740 0.000 40.860 1.120 ;
  LAYER metal4 ;
  RECT 39.740 0.000 40.860 1.120 ;
  LAYER metal3 ;
  RECT 39.740 0.000 40.860 1.120 ;
  LAYER metal2 ;
  RECT 39.740 0.000 40.860 1.120 ;
  LAYER metal1 ;
  RECT 39.740 0.000 40.860 1.120 ;
 END
END DOA1
PIN DIA0
  DIRECTION INPUT ;
  CAPACITANCE 0.010 ;
 PORT
  LAYER metal5 ;
  RECT 26.100 0.000 27.220 1.120 ;
  LAYER metal4 ;
  RECT 26.100 0.000 27.220 1.120 ;
  LAYER metal3 ;
  RECT 26.100 0.000 27.220 1.120 ;
  LAYER metal2 ;
  RECT 26.100 0.000 27.220 1.120 ;
  LAYER metal1 ;
  RECT 26.100 0.000 27.220 1.120 ;
 END
END DIA0
PIN DOA0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.028 ;
 PORT
  LAYER metal5 ;
  RECT 12.460 0.000 13.580 1.120 ;
  LAYER metal4 ;
  RECT 12.460 0.000 13.580 1.120 ;
  LAYER metal3 ;
  RECT 12.460 0.000 13.580 1.120 ;
  LAYER metal2 ;
  RECT 12.460 0.000 13.580 1.120 ;
  LAYER metal1 ;
  RECT 12.460 0.000 13.580 1.120 ;
 END
END DOA0
OBS
  LAYER metal1 SPACING 0.280 ;
  RECT 0.000 0.140 3571.820 209.860 ;
  LAYER metal2 SPACING 0.320 ;
  RECT 0.000 0.140 3571.820 209.860 ;
  LAYER metal3 SPACING 0.320 ;
  RECT 0.000 0.140 3571.820 209.860 ;
  LAYER metal4 SPACING 0.600 ;
  RECT 0.000 0.140 3571.820 209.860 ;
  LAYER via ;
  RECT 0.000 0.140 3571.820 209.860 ;
  LAYER via2 ;
  RECT 0.000 0.140 3571.820 209.860 ;
  LAYER via3 ;
  RECT 0.000 0.140 3571.820 209.860 ;
END
END layer4_sram
END LIBRARY



