# 
#              Synchronous High Speed Single Port SRAM Compiler 
# 
#                    UMC 0.18um GenericII Logic Process
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2009 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http://www.faraday-tech.com/
#   
#       Module Name      : dma_sram
#       Words            : 3072
#       Bits             : 32
#       Byte-Write       : 1
#       Aspect Ratio     : 1
#       Output Loading   : 0.5  (pf)
#       Data Slew        : 2.0  (ns)
#       CK Slew          : 2.0  (ns)
#       Power Ring Width : 2  (um)
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSA0M_A
#       Memaker          : 200901.2.1
#       Date             : 2021/01/15 13:32:42
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO dma_sram
CLASS BLOCK ;
FOREIGN dma_sram 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 563.580 BY 1078.000 ;
SYMMETRY x y r90 ;
SITE core ;
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal4 ;
  RECT 562.460 1066.580 563.580 1069.820 ;
  LAYER metal3 ;
  RECT 562.460 1066.580 563.580 1069.820 ;
  LAYER metal2 ;
  RECT 562.460 1066.580 563.580 1069.820 ;
  LAYER metal1 ;
  RECT 562.460 1066.580 563.580 1069.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 1058.740 563.580 1061.980 ;
  LAYER metal3 ;
  RECT 562.460 1058.740 563.580 1061.980 ;
  LAYER metal2 ;
  RECT 562.460 1058.740 563.580 1061.980 ;
  LAYER metal1 ;
  RECT 562.460 1058.740 563.580 1061.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 1050.900 563.580 1054.140 ;
  LAYER metal3 ;
  RECT 562.460 1050.900 563.580 1054.140 ;
  LAYER metal2 ;
  RECT 562.460 1050.900 563.580 1054.140 ;
  LAYER metal1 ;
  RECT 562.460 1050.900 563.580 1054.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 1043.060 563.580 1046.300 ;
  LAYER metal3 ;
  RECT 562.460 1043.060 563.580 1046.300 ;
  LAYER metal2 ;
  RECT 562.460 1043.060 563.580 1046.300 ;
  LAYER metal1 ;
  RECT 562.460 1043.060 563.580 1046.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 1035.220 563.580 1038.460 ;
  LAYER metal3 ;
  RECT 562.460 1035.220 563.580 1038.460 ;
  LAYER metal2 ;
  RECT 562.460 1035.220 563.580 1038.460 ;
  LAYER metal1 ;
  RECT 562.460 1035.220 563.580 1038.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 1027.380 563.580 1030.620 ;
  LAYER metal3 ;
  RECT 562.460 1027.380 563.580 1030.620 ;
  LAYER metal2 ;
  RECT 562.460 1027.380 563.580 1030.620 ;
  LAYER metal1 ;
  RECT 562.460 1027.380 563.580 1030.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 988.180 563.580 991.420 ;
  LAYER metal3 ;
  RECT 562.460 988.180 563.580 991.420 ;
  LAYER metal2 ;
  RECT 562.460 988.180 563.580 991.420 ;
  LAYER metal1 ;
  RECT 562.460 988.180 563.580 991.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 980.340 563.580 983.580 ;
  LAYER metal3 ;
  RECT 562.460 980.340 563.580 983.580 ;
  LAYER metal2 ;
  RECT 562.460 980.340 563.580 983.580 ;
  LAYER metal1 ;
  RECT 562.460 980.340 563.580 983.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 972.500 563.580 975.740 ;
  LAYER metal3 ;
  RECT 562.460 972.500 563.580 975.740 ;
  LAYER metal2 ;
  RECT 562.460 972.500 563.580 975.740 ;
  LAYER metal1 ;
  RECT 562.460 972.500 563.580 975.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 964.660 563.580 967.900 ;
  LAYER metal3 ;
  RECT 562.460 964.660 563.580 967.900 ;
  LAYER metal2 ;
  RECT 562.460 964.660 563.580 967.900 ;
  LAYER metal1 ;
  RECT 562.460 964.660 563.580 967.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 956.820 563.580 960.060 ;
  LAYER metal3 ;
  RECT 562.460 956.820 563.580 960.060 ;
  LAYER metal2 ;
  RECT 562.460 956.820 563.580 960.060 ;
  LAYER metal1 ;
  RECT 562.460 956.820 563.580 960.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 948.980 563.580 952.220 ;
  LAYER metal3 ;
  RECT 562.460 948.980 563.580 952.220 ;
  LAYER metal2 ;
  RECT 562.460 948.980 563.580 952.220 ;
  LAYER metal1 ;
  RECT 562.460 948.980 563.580 952.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 909.780 563.580 913.020 ;
  LAYER metal3 ;
  RECT 562.460 909.780 563.580 913.020 ;
  LAYER metal2 ;
  RECT 562.460 909.780 563.580 913.020 ;
  LAYER metal1 ;
  RECT 562.460 909.780 563.580 913.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 901.940 563.580 905.180 ;
  LAYER metal3 ;
  RECT 562.460 901.940 563.580 905.180 ;
  LAYER metal2 ;
  RECT 562.460 901.940 563.580 905.180 ;
  LAYER metal1 ;
  RECT 562.460 901.940 563.580 905.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 894.100 563.580 897.340 ;
  LAYER metal3 ;
  RECT 562.460 894.100 563.580 897.340 ;
  LAYER metal2 ;
  RECT 562.460 894.100 563.580 897.340 ;
  LAYER metal1 ;
  RECT 562.460 894.100 563.580 897.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 886.260 563.580 889.500 ;
  LAYER metal3 ;
  RECT 562.460 886.260 563.580 889.500 ;
  LAYER metal2 ;
  RECT 562.460 886.260 563.580 889.500 ;
  LAYER metal1 ;
  RECT 562.460 886.260 563.580 889.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 878.420 563.580 881.660 ;
  LAYER metal3 ;
  RECT 562.460 878.420 563.580 881.660 ;
  LAYER metal2 ;
  RECT 562.460 878.420 563.580 881.660 ;
  LAYER metal1 ;
  RECT 562.460 878.420 563.580 881.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 870.580 563.580 873.820 ;
  LAYER metal3 ;
  RECT 562.460 870.580 563.580 873.820 ;
  LAYER metal2 ;
  RECT 562.460 870.580 563.580 873.820 ;
  LAYER metal1 ;
  RECT 562.460 870.580 563.580 873.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 831.380 563.580 834.620 ;
  LAYER metal3 ;
  RECT 562.460 831.380 563.580 834.620 ;
  LAYER metal2 ;
  RECT 562.460 831.380 563.580 834.620 ;
  LAYER metal1 ;
  RECT 562.460 831.380 563.580 834.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 823.540 563.580 826.780 ;
  LAYER metal3 ;
  RECT 562.460 823.540 563.580 826.780 ;
  LAYER metal2 ;
  RECT 562.460 823.540 563.580 826.780 ;
  LAYER metal1 ;
  RECT 562.460 823.540 563.580 826.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 815.700 563.580 818.940 ;
  LAYER metal3 ;
  RECT 562.460 815.700 563.580 818.940 ;
  LAYER metal2 ;
  RECT 562.460 815.700 563.580 818.940 ;
  LAYER metal1 ;
  RECT 562.460 815.700 563.580 818.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 807.860 563.580 811.100 ;
  LAYER metal3 ;
  RECT 562.460 807.860 563.580 811.100 ;
  LAYER metal2 ;
  RECT 562.460 807.860 563.580 811.100 ;
  LAYER metal1 ;
  RECT 562.460 807.860 563.580 811.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 800.020 563.580 803.260 ;
  LAYER metal3 ;
  RECT 562.460 800.020 563.580 803.260 ;
  LAYER metal2 ;
  RECT 562.460 800.020 563.580 803.260 ;
  LAYER metal1 ;
  RECT 562.460 800.020 563.580 803.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 792.180 563.580 795.420 ;
  LAYER metal3 ;
  RECT 562.460 792.180 563.580 795.420 ;
  LAYER metal2 ;
  RECT 562.460 792.180 563.580 795.420 ;
  LAYER metal1 ;
  RECT 562.460 792.180 563.580 795.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 752.980 563.580 756.220 ;
  LAYER metal3 ;
  RECT 562.460 752.980 563.580 756.220 ;
  LAYER metal2 ;
  RECT 562.460 752.980 563.580 756.220 ;
  LAYER metal1 ;
  RECT 562.460 752.980 563.580 756.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 745.140 563.580 748.380 ;
  LAYER metal3 ;
  RECT 562.460 745.140 563.580 748.380 ;
  LAYER metal2 ;
  RECT 562.460 745.140 563.580 748.380 ;
  LAYER metal1 ;
  RECT 562.460 745.140 563.580 748.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 737.300 563.580 740.540 ;
  LAYER metal3 ;
  RECT 562.460 737.300 563.580 740.540 ;
  LAYER metal2 ;
  RECT 562.460 737.300 563.580 740.540 ;
  LAYER metal1 ;
  RECT 562.460 737.300 563.580 740.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 729.460 563.580 732.700 ;
  LAYER metal3 ;
  RECT 562.460 729.460 563.580 732.700 ;
  LAYER metal2 ;
  RECT 562.460 729.460 563.580 732.700 ;
  LAYER metal1 ;
  RECT 562.460 729.460 563.580 732.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 721.620 563.580 724.860 ;
  LAYER metal3 ;
  RECT 562.460 721.620 563.580 724.860 ;
  LAYER metal2 ;
  RECT 562.460 721.620 563.580 724.860 ;
  LAYER metal1 ;
  RECT 562.460 721.620 563.580 724.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 713.780 563.580 717.020 ;
  LAYER metal3 ;
  RECT 562.460 713.780 563.580 717.020 ;
  LAYER metal2 ;
  RECT 562.460 713.780 563.580 717.020 ;
  LAYER metal1 ;
  RECT 562.460 713.780 563.580 717.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 674.580 563.580 677.820 ;
  LAYER metal3 ;
  RECT 562.460 674.580 563.580 677.820 ;
  LAYER metal2 ;
  RECT 562.460 674.580 563.580 677.820 ;
  LAYER metal1 ;
  RECT 562.460 674.580 563.580 677.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 666.740 563.580 669.980 ;
  LAYER metal3 ;
  RECT 562.460 666.740 563.580 669.980 ;
  LAYER metal2 ;
  RECT 562.460 666.740 563.580 669.980 ;
  LAYER metal1 ;
  RECT 562.460 666.740 563.580 669.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 658.900 563.580 662.140 ;
  LAYER metal3 ;
  RECT 562.460 658.900 563.580 662.140 ;
  LAYER metal2 ;
  RECT 562.460 658.900 563.580 662.140 ;
  LAYER metal1 ;
  RECT 562.460 658.900 563.580 662.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 651.060 563.580 654.300 ;
  LAYER metal3 ;
  RECT 562.460 651.060 563.580 654.300 ;
  LAYER metal2 ;
  RECT 562.460 651.060 563.580 654.300 ;
  LAYER metal1 ;
  RECT 562.460 651.060 563.580 654.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 643.220 563.580 646.460 ;
  LAYER metal3 ;
  RECT 562.460 643.220 563.580 646.460 ;
  LAYER metal2 ;
  RECT 562.460 643.220 563.580 646.460 ;
  LAYER metal1 ;
  RECT 562.460 643.220 563.580 646.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 635.380 563.580 638.620 ;
  LAYER metal3 ;
  RECT 562.460 635.380 563.580 638.620 ;
  LAYER metal2 ;
  RECT 562.460 635.380 563.580 638.620 ;
  LAYER metal1 ;
  RECT 562.460 635.380 563.580 638.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 596.180 563.580 599.420 ;
  LAYER metal3 ;
  RECT 562.460 596.180 563.580 599.420 ;
  LAYER metal2 ;
  RECT 562.460 596.180 563.580 599.420 ;
  LAYER metal1 ;
  RECT 562.460 596.180 563.580 599.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 588.340 563.580 591.580 ;
  LAYER metal3 ;
  RECT 562.460 588.340 563.580 591.580 ;
  LAYER metal2 ;
  RECT 562.460 588.340 563.580 591.580 ;
  LAYER metal1 ;
  RECT 562.460 588.340 563.580 591.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 580.500 563.580 583.740 ;
  LAYER metal3 ;
  RECT 562.460 580.500 563.580 583.740 ;
  LAYER metal2 ;
  RECT 562.460 580.500 563.580 583.740 ;
  LAYER metal1 ;
  RECT 562.460 580.500 563.580 583.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 572.660 563.580 575.900 ;
  LAYER metal3 ;
  RECT 562.460 572.660 563.580 575.900 ;
  LAYER metal2 ;
  RECT 562.460 572.660 563.580 575.900 ;
  LAYER metal1 ;
  RECT 562.460 572.660 563.580 575.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 564.820 563.580 568.060 ;
  LAYER metal3 ;
  RECT 562.460 564.820 563.580 568.060 ;
  LAYER metal2 ;
  RECT 562.460 564.820 563.580 568.060 ;
  LAYER metal1 ;
  RECT 562.460 564.820 563.580 568.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 556.980 563.580 560.220 ;
  LAYER metal3 ;
  RECT 562.460 556.980 563.580 560.220 ;
  LAYER metal2 ;
  RECT 562.460 556.980 563.580 560.220 ;
  LAYER metal1 ;
  RECT 562.460 556.980 563.580 560.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 517.780 563.580 521.020 ;
  LAYER metal3 ;
  RECT 562.460 517.780 563.580 521.020 ;
  LAYER metal2 ;
  RECT 562.460 517.780 563.580 521.020 ;
  LAYER metal1 ;
  RECT 562.460 517.780 563.580 521.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 509.940 563.580 513.180 ;
  LAYER metal3 ;
  RECT 562.460 509.940 563.580 513.180 ;
  LAYER metal2 ;
  RECT 562.460 509.940 563.580 513.180 ;
  LAYER metal1 ;
  RECT 562.460 509.940 563.580 513.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 502.100 563.580 505.340 ;
  LAYER metal3 ;
  RECT 562.460 502.100 563.580 505.340 ;
  LAYER metal2 ;
  RECT 562.460 502.100 563.580 505.340 ;
  LAYER metal1 ;
  RECT 562.460 502.100 563.580 505.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 494.260 563.580 497.500 ;
  LAYER metal3 ;
  RECT 562.460 494.260 563.580 497.500 ;
  LAYER metal2 ;
  RECT 562.460 494.260 563.580 497.500 ;
  LAYER metal1 ;
  RECT 562.460 494.260 563.580 497.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 486.420 563.580 489.660 ;
  LAYER metal3 ;
  RECT 562.460 486.420 563.580 489.660 ;
  LAYER metal2 ;
  RECT 562.460 486.420 563.580 489.660 ;
  LAYER metal1 ;
  RECT 562.460 486.420 563.580 489.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 478.580 563.580 481.820 ;
  LAYER metal3 ;
  RECT 562.460 478.580 563.580 481.820 ;
  LAYER metal2 ;
  RECT 562.460 478.580 563.580 481.820 ;
  LAYER metal1 ;
  RECT 562.460 478.580 563.580 481.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 439.380 563.580 442.620 ;
  LAYER metal3 ;
  RECT 562.460 439.380 563.580 442.620 ;
  LAYER metal2 ;
  RECT 562.460 439.380 563.580 442.620 ;
  LAYER metal1 ;
  RECT 562.460 439.380 563.580 442.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 431.540 563.580 434.780 ;
  LAYER metal3 ;
  RECT 562.460 431.540 563.580 434.780 ;
  LAYER metal2 ;
  RECT 562.460 431.540 563.580 434.780 ;
  LAYER metal1 ;
  RECT 562.460 431.540 563.580 434.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 423.700 563.580 426.940 ;
  LAYER metal3 ;
  RECT 562.460 423.700 563.580 426.940 ;
  LAYER metal2 ;
  RECT 562.460 423.700 563.580 426.940 ;
  LAYER metal1 ;
  RECT 562.460 423.700 563.580 426.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 415.860 563.580 419.100 ;
  LAYER metal3 ;
  RECT 562.460 415.860 563.580 419.100 ;
  LAYER metal2 ;
  RECT 562.460 415.860 563.580 419.100 ;
  LAYER metal1 ;
  RECT 562.460 415.860 563.580 419.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 408.020 563.580 411.260 ;
  LAYER metal3 ;
  RECT 562.460 408.020 563.580 411.260 ;
  LAYER metal2 ;
  RECT 562.460 408.020 563.580 411.260 ;
  LAYER metal1 ;
  RECT 562.460 408.020 563.580 411.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 400.180 563.580 403.420 ;
  LAYER metal3 ;
  RECT 562.460 400.180 563.580 403.420 ;
  LAYER metal2 ;
  RECT 562.460 400.180 563.580 403.420 ;
  LAYER metal1 ;
  RECT 562.460 400.180 563.580 403.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 360.980 563.580 364.220 ;
  LAYER metal3 ;
  RECT 562.460 360.980 563.580 364.220 ;
  LAYER metal2 ;
  RECT 562.460 360.980 563.580 364.220 ;
  LAYER metal1 ;
  RECT 562.460 360.980 563.580 364.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 353.140 563.580 356.380 ;
  LAYER metal3 ;
  RECT 562.460 353.140 563.580 356.380 ;
  LAYER metal2 ;
  RECT 562.460 353.140 563.580 356.380 ;
  LAYER metal1 ;
  RECT 562.460 353.140 563.580 356.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 345.300 563.580 348.540 ;
  LAYER metal3 ;
  RECT 562.460 345.300 563.580 348.540 ;
  LAYER metal2 ;
  RECT 562.460 345.300 563.580 348.540 ;
  LAYER metal1 ;
  RECT 562.460 345.300 563.580 348.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 337.460 563.580 340.700 ;
  LAYER metal3 ;
  RECT 562.460 337.460 563.580 340.700 ;
  LAYER metal2 ;
  RECT 562.460 337.460 563.580 340.700 ;
  LAYER metal1 ;
  RECT 562.460 337.460 563.580 340.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 329.620 563.580 332.860 ;
  LAYER metal3 ;
  RECT 562.460 329.620 563.580 332.860 ;
  LAYER metal2 ;
  RECT 562.460 329.620 563.580 332.860 ;
  LAYER metal1 ;
  RECT 562.460 329.620 563.580 332.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 321.780 563.580 325.020 ;
  LAYER metal3 ;
  RECT 562.460 321.780 563.580 325.020 ;
  LAYER metal2 ;
  RECT 562.460 321.780 563.580 325.020 ;
  LAYER metal1 ;
  RECT 562.460 321.780 563.580 325.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 282.580 563.580 285.820 ;
  LAYER metal3 ;
  RECT 562.460 282.580 563.580 285.820 ;
  LAYER metal2 ;
  RECT 562.460 282.580 563.580 285.820 ;
  LAYER metal1 ;
  RECT 562.460 282.580 563.580 285.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 274.740 563.580 277.980 ;
  LAYER metal3 ;
  RECT 562.460 274.740 563.580 277.980 ;
  LAYER metal2 ;
  RECT 562.460 274.740 563.580 277.980 ;
  LAYER metal1 ;
  RECT 562.460 274.740 563.580 277.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 266.900 563.580 270.140 ;
  LAYER metal3 ;
  RECT 562.460 266.900 563.580 270.140 ;
  LAYER metal2 ;
  RECT 562.460 266.900 563.580 270.140 ;
  LAYER metal1 ;
  RECT 562.460 266.900 563.580 270.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 259.060 563.580 262.300 ;
  LAYER metal3 ;
  RECT 562.460 259.060 563.580 262.300 ;
  LAYER metal2 ;
  RECT 562.460 259.060 563.580 262.300 ;
  LAYER metal1 ;
  RECT 562.460 259.060 563.580 262.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 251.220 563.580 254.460 ;
  LAYER metal3 ;
  RECT 562.460 251.220 563.580 254.460 ;
  LAYER metal2 ;
  RECT 562.460 251.220 563.580 254.460 ;
  LAYER metal1 ;
  RECT 562.460 251.220 563.580 254.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 243.380 563.580 246.620 ;
  LAYER metal3 ;
  RECT 562.460 243.380 563.580 246.620 ;
  LAYER metal2 ;
  RECT 562.460 243.380 563.580 246.620 ;
  LAYER metal1 ;
  RECT 562.460 243.380 563.580 246.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 204.180 563.580 207.420 ;
  LAYER metal3 ;
  RECT 562.460 204.180 563.580 207.420 ;
  LAYER metal2 ;
  RECT 562.460 204.180 563.580 207.420 ;
  LAYER metal1 ;
  RECT 562.460 204.180 563.580 207.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 196.340 563.580 199.580 ;
  LAYER metal3 ;
  RECT 562.460 196.340 563.580 199.580 ;
  LAYER metal2 ;
  RECT 562.460 196.340 563.580 199.580 ;
  LAYER metal1 ;
  RECT 562.460 196.340 563.580 199.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 188.500 563.580 191.740 ;
  LAYER metal3 ;
  RECT 562.460 188.500 563.580 191.740 ;
  LAYER metal2 ;
  RECT 562.460 188.500 563.580 191.740 ;
  LAYER metal1 ;
  RECT 562.460 188.500 563.580 191.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 180.660 563.580 183.900 ;
  LAYER metal3 ;
  RECT 562.460 180.660 563.580 183.900 ;
  LAYER metal2 ;
  RECT 562.460 180.660 563.580 183.900 ;
  LAYER metal1 ;
  RECT 562.460 180.660 563.580 183.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 172.820 563.580 176.060 ;
  LAYER metal3 ;
  RECT 562.460 172.820 563.580 176.060 ;
  LAYER metal2 ;
  RECT 562.460 172.820 563.580 176.060 ;
  LAYER metal1 ;
  RECT 562.460 172.820 563.580 176.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 164.980 563.580 168.220 ;
  LAYER metal3 ;
  RECT 562.460 164.980 563.580 168.220 ;
  LAYER metal2 ;
  RECT 562.460 164.980 563.580 168.220 ;
  LAYER metal1 ;
  RECT 562.460 164.980 563.580 168.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 125.780 563.580 129.020 ;
  LAYER metal3 ;
  RECT 562.460 125.780 563.580 129.020 ;
  LAYER metal2 ;
  RECT 562.460 125.780 563.580 129.020 ;
  LAYER metal1 ;
  RECT 562.460 125.780 563.580 129.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 117.940 563.580 121.180 ;
  LAYER metal3 ;
  RECT 562.460 117.940 563.580 121.180 ;
  LAYER metal2 ;
  RECT 562.460 117.940 563.580 121.180 ;
  LAYER metal1 ;
  RECT 562.460 117.940 563.580 121.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 110.100 563.580 113.340 ;
  LAYER metal3 ;
  RECT 562.460 110.100 563.580 113.340 ;
  LAYER metal2 ;
  RECT 562.460 110.100 563.580 113.340 ;
  LAYER metal1 ;
  RECT 562.460 110.100 563.580 113.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 102.260 563.580 105.500 ;
  LAYER metal3 ;
  RECT 562.460 102.260 563.580 105.500 ;
  LAYER metal2 ;
  RECT 562.460 102.260 563.580 105.500 ;
  LAYER metal1 ;
  RECT 562.460 102.260 563.580 105.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 94.420 563.580 97.660 ;
  LAYER metal3 ;
  RECT 562.460 94.420 563.580 97.660 ;
  LAYER metal2 ;
  RECT 562.460 94.420 563.580 97.660 ;
  LAYER metal1 ;
  RECT 562.460 94.420 563.580 97.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 86.580 563.580 89.820 ;
  LAYER metal3 ;
  RECT 562.460 86.580 563.580 89.820 ;
  LAYER metal2 ;
  RECT 562.460 86.580 563.580 89.820 ;
  LAYER metal1 ;
  RECT 562.460 86.580 563.580 89.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 47.380 563.580 50.620 ;
  LAYER metal3 ;
  RECT 562.460 47.380 563.580 50.620 ;
  LAYER metal2 ;
  RECT 562.460 47.380 563.580 50.620 ;
  LAYER metal1 ;
  RECT 562.460 47.380 563.580 50.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 39.540 563.580 42.780 ;
  LAYER metal3 ;
  RECT 562.460 39.540 563.580 42.780 ;
  LAYER metal2 ;
  RECT 562.460 39.540 563.580 42.780 ;
  LAYER metal1 ;
  RECT 562.460 39.540 563.580 42.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 31.700 563.580 34.940 ;
  LAYER metal3 ;
  RECT 562.460 31.700 563.580 34.940 ;
  LAYER metal2 ;
  RECT 562.460 31.700 563.580 34.940 ;
  LAYER metal1 ;
  RECT 562.460 31.700 563.580 34.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 23.860 563.580 27.100 ;
  LAYER metal3 ;
  RECT 562.460 23.860 563.580 27.100 ;
  LAYER metal2 ;
  RECT 562.460 23.860 563.580 27.100 ;
  LAYER metal1 ;
  RECT 562.460 23.860 563.580 27.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 16.020 563.580 19.260 ;
  LAYER metal3 ;
  RECT 562.460 16.020 563.580 19.260 ;
  LAYER metal2 ;
  RECT 562.460 16.020 563.580 19.260 ;
  LAYER metal1 ;
  RECT 562.460 16.020 563.580 19.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 8.180 563.580 11.420 ;
  LAYER metal3 ;
  RECT 562.460 8.180 563.580 11.420 ;
  LAYER metal2 ;
  RECT 562.460 8.180 563.580 11.420 ;
  LAYER metal1 ;
  RECT 562.460 8.180 563.580 11.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1066.580 1.120 1069.820 ;
  LAYER metal3 ;
  RECT 0.000 1066.580 1.120 1069.820 ;
  LAYER metal2 ;
  RECT 0.000 1066.580 1.120 1069.820 ;
  LAYER metal1 ;
  RECT 0.000 1066.580 1.120 1069.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1058.740 1.120 1061.980 ;
  LAYER metal3 ;
  RECT 0.000 1058.740 1.120 1061.980 ;
  LAYER metal2 ;
  RECT 0.000 1058.740 1.120 1061.980 ;
  LAYER metal1 ;
  RECT 0.000 1058.740 1.120 1061.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1050.900 1.120 1054.140 ;
  LAYER metal3 ;
  RECT 0.000 1050.900 1.120 1054.140 ;
  LAYER metal2 ;
  RECT 0.000 1050.900 1.120 1054.140 ;
  LAYER metal1 ;
  RECT 0.000 1050.900 1.120 1054.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1043.060 1.120 1046.300 ;
  LAYER metal3 ;
  RECT 0.000 1043.060 1.120 1046.300 ;
  LAYER metal2 ;
  RECT 0.000 1043.060 1.120 1046.300 ;
  LAYER metal1 ;
  RECT 0.000 1043.060 1.120 1046.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1035.220 1.120 1038.460 ;
  LAYER metal3 ;
  RECT 0.000 1035.220 1.120 1038.460 ;
  LAYER metal2 ;
  RECT 0.000 1035.220 1.120 1038.460 ;
  LAYER metal1 ;
  RECT 0.000 1035.220 1.120 1038.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1027.380 1.120 1030.620 ;
  LAYER metal3 ;
  RECT 0.000 1027.380 1.120 1030.620 ;
  LAYER metal2 ;
  RECT 0.000 1027.380 1.120 1030.620 ;
  LAYER metal1 ;
  RECT 0.000 1027.380 1.120 1030.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 988.180 1.120 991.420 ;
  LAYER metal3 ;
  RECT 0.000 988.180 1.120 991.420 ;
  LAYER metal2 ;
  RECT 0.000 988.180 1.120 991.420 ;
  LAYER metal1 ;
  RECT 0.000 988.180 1.120 991.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 980.340 1.120 983.580 ;
  LAYER metal3 ;
  RECT 0.000 980.340 1.120 983.580 ;
  LAYER metal2 ;
  RECT 0.000 980.340 1.120 983.580 ;
  LAYER metal1 ;
  RECT 0.000 980.340 1.120 983.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 972.500 1.120 975.740 ;
  LAYER metal3 ;
  RECT 0.000 972.500 1.120 975.740 ;
  LAYER metal2 ;
  RECT 0.000 972.500 1.120 975.740 ;
  LAYER metal1 ;
  RECT 0.000 972.500 1.120 975.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 964.660 1.120 967.900 ;
  LAYER metal3 ;
  RECT 0.000 964.660 1.120 967.900 ;
  LAYER metal2 ;
  RECT 0.000 964.660 1.120 967.900 ;
  LAYER metal1 ;
  RECT 0.000 964.660 1.120 967.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 956.820 1.120 960.060 ;
  LAYER metal3 ;
  RECT 0.000 956.820 1.120 960.060 ;
  LAYER metal2 ;
  RECT 0.000 956.820 1.120 960.060 ;
  LAYER metal1 ;
  RECT 0.000 956.820 1.120 960.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 948.980 1.120 952.220 ;
  LAYER metal3 ;
  RECT 0.000 948.980 1.120 952.220 ;
  LAYER metal2 ;
  RECT 0.000 948.980 1.120 952.220 ;
  LAYER metal1 ;
  RECT 0.000 948.980 1.120 952.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 909.780 1.120 913.020 ;
  LAYER metal3 ;
  RECT 0.000 909.780 1.120 913.020 ;
  LAYER metal2 ;
  RECT 0.000 909.780 1.120 913.020 ;
  LAYER metal1 ;
  RECT 0.000 909.780 1.120 913.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 901.940 1.120 905.180 ;
  LAYER metal3 ;
  RECT 0.000 901.940 1.120 905.180 ;
  LAYER metal2 ;
  RECT 0.000 901.940 1.120 905.180 ;
  LAYER metal1 ;
  RECT 0.000 901.940 1.120 905.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 894.100 1.120 897.340 ;
  LAYER metal3 ;
  RECT 0.000 894.100 1.120 897.340 ;
  LAYER metal2 ;
  RECT 0.000 894.100 1.120 897.340 ;
  LAYER metal1 ;
  RECT 0.000 894.100 1.120 897.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 886.260 1.120 889.500 ;
  LAYER metal3 ;
  RECT 0.000 886.260 1.120 889.500 ;
  LAYER metal2 ;
  RECT 0.000 886.260 1.120 889.500 ;
  LAYER metal1 ;
  RECT 0.000 886.260 1.120 889.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 878.420 1.120 881.660 ;
  LAYER metal3 ;
  RECT 0.000 878.420 1.120 881.660 ;
  LAYER metal2 ;
  RECT 0.000 878.420 1.120 881.660 ;
  LAYER metal1 ;
  RECT 0.000 878.420 1.120 881.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 870.580 1.120 873.820 ;
  LAYER metal3 ;
  RECT 0.000 870.580 1.120 873.820 ;
  LAYER metal2 ;
  RECT 0.000 870.580 1.120 873.820 ;
  LAYER metal1 ;
  RECT 0.000 870.580 1.120 873.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 831.380 1.120 834.620 ;
  LAYER metal3 ;
  RECT 0.000 831.380 1.120 834.620 ;
  LAYER metal2 ;
  RECT 0.000 831.380 1.120 834.620 ;
  LAYER metal1 ;
  RECT 0.000 831.380 1.120 834.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 823.540 1.120 826.780 ;
  LAYER metal3 ;
  RECT 0.000 823.540 1.120 826.780 ;
  LAYER metal2 ;
  RECT 0.000 823.540 1.120 826.780 ;
  LAYER metal1 ;
  RECT 0.000 823.540 1.120 826.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 815.700 1.120 818.940 ;
  LAYER metal3 ;
  RECT 0.000 815.700 1.120 818.940 ;
  LAYER metal2 ;
  RECT 0.000 815.700 1.120 818.940 ;
  LAYER metal1 ;
  RECT 0.000 815.700 1.120 818.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 807.860 1.120 811.100 ;
  LAYER metal3 ;
  RECT 0.000 807.860 1.120 811.100 ;
  LAYER metal2 ;
  RECT 0.000 807.860 1.120 811.100 ;
  LAYER metal1 ;
  RECT 0.000 807.860 1.120 811.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 800.020 1.120 803.260 ;
  LAYER metal3 ;
  RECT 0.000 800.020 1.120 803.260 ;
  LAYER metal2 ;
  RECT 0.000 800.020 1.120 803.260 ;
  LAYER metal1 ;
  RECT 0.000 800.020 1.120 803.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 792.180 1.120 795.420 ;
  LAYER metal3 ;
  RECT 0.000 792.180 1.120 795.420 ;
  LAYER metal2 ;
  RECT 0.000 792.180 1.120 795.420 ;
  LAYER metal1 ;
  RECT 0.000 792.180 1.120 795.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 752.980 1.120 756.220 ;
  LAYER metal3 ;
  RECT 0.000 752.980 1.120 756.220 ;
  LAYER metal2 ;
  RECT 0.000 752.980 1.120 756.220 ;
  LAYER metal1 ;
  RECT 0.000 752.980 1.120 756.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 745.140 1.120 748.380 ;
  LAYER metal3 ;
  RECT 0.000 745.140 1.120 748.380 ;
  LAYER metal2 ;
  RECT 0.000 745.140 1.120 748.380 ;
  LAYER metal1 ;
  RECT 0.000 745.140 1.120 748.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 737.300 1.120 740.540 ;
  LAYER metal3 ;
  RECT 0.000 737.300 1.120 740.540 ;
  LAYER metal2 ;
  RECT 0.000 737.300 1.120 740.540 ;
  LAYER metal1 ;
  RECT 0.000 737.300 1.120 740.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 729.460 1.120 732.700 ;
  LAYER metal3 ;
  RECT 0.000 729.460 1.120 732.700 ;
  LAYER metal2 ;
  RECT 0.000 729.460 1.120 732.700 ;
  LAYER metal1 ;
  RECT 0.000 729.460 1.120 732.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 721.620 1.120 724.860 ;
  LAYER metal3 ;
  RECT 0.000 721.620 1.120 724.860 ;
  LAYER metal2 ;
  RECT 0.000 721.620 1.120 724.860 ;
  LAYER metal1 ;
  RECT 0.000 721.620 1.120 724.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 713.780 1.120 717.020 ;
  LAYER metal3 ;
  RECT 0.000 713.780 1.120 717.020 ;
  LAYER metal2 ;
  RECT 0.000 713.780 1.120 717.020 ;
  LAYER metal1 ;
  RECT 0.000 713.780 1.120 717.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 674.580 1.120 677.820 ;
  LAYER metal3 ;
  RECT 0.000 674.580 1.120 677.820 ;
  LAYER metal2 ;
  RECT 0.000 674.580 1.120 677.820 ;
  LAYER metal1 ;
  RECT 0.000 674.580 1.120 677.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 666.740 1.120 669.980 ;
  LAYER metal3 ;
  RECT 0.000 666.740 1.120 669.980 ;
  LAYER metal2 ;
  RECT 0.000 666.740 1.120 669.980 ;
  LAYER metal1 ;
  RECT 0.000 666.740 1.120 669.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 658.900 1.120 662.140 ;
  LAYER metal3 ;
  RECT 0.000 658.900 1.120 662.140 ;
  LAYER metal2 ;
  RECT 0.000 658.900 1.120 662.140 ;
  LAYER metal1 ;
  RECT 0.000 658.900 1.120 662.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 651.060 1.120 654.300 ;
  LAYER metal3 ;
  RECT 0.000 651.060 1.120 654.300 ;
  LAYER metal2 ;
  RECT 0.000 651.060 1.120 654.300 ;
  LAYER metal1 ;
  RECT 0.000 651.060 1.120 654.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 643.220 1.120 646.460 ;
  LAYER metal3 ;
  RECT 0.000 643.220 1.120 646.460 ;
  LAYER metal2 ;
  RECT 0.000 643.220 1.120 646.460 ;
  LAYER metal1 ;
  RECT 0.000 643.220 1.120 646.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 635.380 1.120 638.620 ;
  LAYER metal3 ;
  RECT 0.000 635.380 1.120 638.620 ;
  LAYER metal2 ;
  RECT 0.000 635.380 1.120 638.620 ;
  LAYER metal1 ;
  RECT 0.000 635.380 1.120 638.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 596.180 1.120 599.420 ;
  LAYER metal3 ;
  RECT 0.000 596.180 1.120 599.420 ;
  LAYER metal2 ;
  RECT 0.000 596.180 1.120 599.420 ;
  LAYER metal1 ;
  RECT 0.000 596.180 1.120 599.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 588.340 1.120 591.580 ;
  LAYER metal3 ;
  RECT 0.000 588.340 1.120 591.580 ;
  LAYER metal2 ;
  RECT 0.000 588.340 1.120 591.580 ;
  LAYER metal1 ;
  RECT 0.000 588.340 1.120 591.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 580.500 1.120 583.740 ;
  LAYER metal3 ;
  RECT 0.000 580.500 1.120 583.740 ;
  LAYER metal2 ;
  RECT 0.000 580.500 1.120 583.740 ;
  LAYER metal1 ;
  RECT 0.000 580.500 1.120 583.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 572.660 1.120 575.900 ;
  LAYER metal3 ;
  RECT 0.000 572.660 1.120 575.900 ;
  LAYER metal2 ;
  RECT 0.000 572.660 1.120 575.900 ;
  LAYER metal1 ;
  RECT 0.000 572.660 1.120 575.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 564.820 1.120 568.060 ;
  LAYER metal3 ;
  RECT 0.000 564.820 1.120 568.060 ;
  LAYER metal2 ;
  RECT 0.000 564.820 1.120 568.060 ;
  LAYER metal1 ;
  RECT 0.000 564.820 1.120 568.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 556.980 1.120 560.220 ;
  LAYER metal3 ;
  RECT 0.000 556.980 1.120 560.220 ;
  LAYER metal2 ;
  RECT 0.000 556.980 1.120 560.220 ;
  LAYER metal1 ;
  RECT 0.000 556.980 1.120 560.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 517.780 1.120 521.020 ;
  LAYER metal3 ;
  RECT 0.000 517.780 1.120 521.020 ;
  LAYER metal2 ;
  RECT 0.000 517.780 1.120 521.020 ;
  LAYER metal1 ;
  RECT 0.000 517.780 1.120 521.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 509.940 1.120 513.180 ;
  LAYER metal3 ;
  RECT 0.000 509.940 1.120 513.180 ;
  LAYER metal2 ;
  RECT 0.000 509.940 1.120 513.180 ;
  LAYER metal1 ;
  RECT 0.000 509.940 1.120 513.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 502.100 1.120 505.340 ;
  LAYER metal3 ;
  RECT 0.000 502.100 1.120 505.340 ;
  LAYER metal2 ;
  RECT 0.000 502.100 1.120 505.340 ;
  LAYER metal1 ;
  RECT 0.000 502.100 1.120 505.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 494.260 1.120 497.500 ;
  LAYER metal3 ;
  RECT 0.000 494.260 1.120 497.500 ;
  LAYER metal2 ;
  RECT 0.000 494.260 1.120 497.500 ;
  LAYER metal1 ;
  RECT 0.000 494.260 1.120 497.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 486.420 1.120 489.660 ;
  LAYER metal3 ;
  RECT 0.000 486.420 1.120 489.660 ;
  LAYER metal2 ;
  RECT 0.000 486.420 1.120 489.660 ;
  LAYER metal1 ;
  RECT 0.000 486.420 1.120 489.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 478.580 1.120 481.820 ;
  LAYER metal3 ;
  RECT 0.000 478.580 1.120 481.820 ;
  LAYER metal2 ;
  RECT 0.000 478.580 1.120 481.820 ;
  LAYER metal1 ;
  RECT 0.000 478.580 1.120 481.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 439.380 1.120 442.620 ;
  LAYER metal3 ;
  RECT 0.000 439.380 1.120 442.620 ;
  LAYER metal2 ;
  RECT 0.000 439.380 1.120 442.620 ;
  LAYER metal1 ;
  RECT 0.000 439.380 1.120 442.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 431.540 1.120 434.780 ;
  LAYER metal3 ;
  RECT 0.000 431.540 1.120 434.780 ;
  LAYER metal2 ;
  RECT 0.000 431.540 1.120 434.780 ;
  LAYER metal1 ;
  RECT 0.000 431.540 1.120 434.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 423.700 1.120 426.940 ;
  LAYER metal3 ;
  RECT 0.000 423.700 1.120 426.940 ;
  LAYER metal2 ;
  RECT 0.000 423.700 1.120 426.940 ;
  LAYER metal1 ;
  RECT 0.000 423.700 1.120 426.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 415.860 1.120 419.100 ;
  LAYER metal3 ;
  RECT 0.000 415.860 1.120 419.100 ;
  LAYER metal2 ;
  RECT 0.000 415.860 1.120 419.100 ;
  LAYER metal1 ;
  RECT 0.000 415.860 1.120 419.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 408.020 1.120 411.260 ;
  LAYER metal3 ;
  RECT 0.000 408.020 1.120 411.260 ;
  LAYER metal2 ;
  RECT 0.000 408.020 1.120 411.260 ;
  LAYER metal1 ;
  RECT 0.000 408.020 1.120 411.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 400.180 1.120 403.420 ;
  LAYER metal3 ;
  RECT 0.000 400.180 1.120 403.420 ;
  LAYER metal2 ;
  RECT 0.000 400.180 1.120 403.420 ;
  LAYER metal1 ;
  RECT 0.000 400.180 1.120 403.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 360.980 1.120 364.220 ;
  LAYER metal3 ;
  RECT 0.000 360.980 1.120 364.220 ;
  LAYER metal2 ;
  RECT 0.000 360.980 1.120 364.220 ;
  LAYER metal1 ;
  RECT 0.000 360.980 1.120 364.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 353.140 1.120 356.380 ;
  LAYER metal3 ;
  RECT 0.000 353.140 1.120 356.380 ;
  LAYER metal2 ;
  RECT 0.000 353.140 1.120 356.380 ;
  LAYER metal1 ;
  RECT 0.000 353.140 1.120 356.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 345.300 1.120 348.540 ;
  LAYER metal3 ;
  RECT 0.000 345.300 1.120 348.540 ;
  LAYER metal2 ;
  RECT 0.000 345.300 1.120 348.540 ;
  LAYER metal1 ;
  RECT 0.000 345.300 1.120 348.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 337.460 1.120 340.700 ;
  LAYER metal3 ;
  RECT 0.000 337.460 1.120 340.700 ;
  LAYER metal2 ;
  RECT 0.000 337.460 1.120 340.700 ;
  LAYER metal1 ;
  RECT 0.000 337.460 1.120 340.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 329.620 1.120 332.860 ;
  LAYER metal3 ;
  RECT 0.000 329.620 1.120 332.860 ;
  LAYER metal2 ;
  RECT 0.000 329.620 1.120 332.860 ;
  LAYER metal1 ;
  RECT 0.000 329.620 1.120 332.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 321.780 1.120 325.020 ;
  LAYER metal3 ;
  RECT 0.000 321.780 1.120 325.020 ;
  LAYER metal2 ;
  RECT 0.000 321.780 1.120 325.020 ;
  LAYER metal1 ;
  RECT 0.000 321.780 1.120 325.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 282.580 1.120 285.820 ;
  LAYER metal3 ;
  RECT 0.000 282.580 1.120 285.820 ;
  LAYER metal2 ;
  RECT 0.000 282.580 1.120 285.820 ;
  LAYER metal1 ;
  RECT 0.000 282.580 1.120 285.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 274.740 1.120 277.980 ;
  LAYER metal3 ;
  RECT 0.000 274.740 1.120 277.980 ;
  LAYER metal2 ;
  RECT 0.000 274.740 1.120 277.980 ;
  LAYER metal1 ;
  RECT 0.000 274.740 1.120 277.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 266.900 1.120 270.140 ;
  LAYER metal3 ;
  RECT 0.000 266.900 1.120 270.140 ;
  LAYER metal2 ;
  RECT 0.000 266.900 1.120 270.140 ;
  LAYER metal1 ;
  RECT 0.000 266.900 1.120 270.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 259.060 1.120 262.300 ;
  LAYER metal3 ;
  RECT 0.000 259.060 1.120 262.300 ;
  LAYER metal2 ;
  RECT 0.000 259.060 1.120 262.300 ;
  LAYER metal1 ;
  RECT 0.000 259.060 1.120 262.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 251.220 1.120 254.460 ;
  LAYER metal3 ;
  RECT 0.000 251.220 1.120 254.460 ;
  LAYER metal2 ;
  RECT 0.000 251.220 1.120 254.460 ;
  LAYER metal1 ;
  RECT 0.000 251.220 1.120 254.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER metal3 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER metal2 ;
  RECT 0.000 243.380 1.120 246.620 ;
  LAYER metal1 ;
  RECT 0.000 243.380 1.120 246.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER metal3 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER metal2 ;
  RECT 0.000 204.180 1.120 207.420 ;
  LAYER metal1 ;
  RECT 0.000 204.180 1.120 207.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER metal3 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER metal2 ;
  RECT 0.000 196.340 1.120 199.580 ;
  LAYER metal1 ;
  RECT 0.000 196.340 1.120 199.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER metal3 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER metal2 ;
  RECT 0.000 188.500 1.120 191.740 ;
  LAYER metal1 ;
  RECT 0.000 188.500 1.120 191.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER metal3 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER metal2 ;
  RECT 0.000 180.660 1.120 183.900 ;
  LAYER metal1 ;
  RECT 0.000 180.660 1.120 183.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER metal3 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER metal2 ;
  RECT 0.000 172.820 1.120 176.060 ;
  LAYER metal1 ;
  RECT 0.000 172.820 1.120 176.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER metal3 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER metal2 ;
  RECT 0.000 164.980 1.120 168.220 ;
  LAYER metal1 ;
  RECT 0.000 164.980 1.120 168.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal3 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal2 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER metal1 ;
  RECT 0.000 125.780 1.120 129.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal3 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal2 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER metal1 ;
  RECT 0.000 117.940 1.120 121.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal3 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal2 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER metal1 ;
  RECT 0.000 110.100 1.120 113.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal3 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal2 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER metal1 ;
  RECT 0.000 102.260 1.120 105.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal3 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal2 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER metal1 ;
  RECT 0.000 94.420 1.120 97.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal3 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal2 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER metal1 ;
  RECT 0.000 86.580 1.120 89.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal3 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal2 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER metal1 ;
  RECT 0.000 47.380 1.120 50.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal3 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal2 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER metal1 ;
  RECT 0.000 39.540 1.120 42.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal3 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal2 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER metal1 ;
  RECT 0.000 31.700 1.120 34.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal3 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal2 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER metal1 ;
  RECT 0.000 23.860 1.120 27.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal3 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal2 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER metal1 ;
  RECT 0.000 16.020 1.120 19.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal3 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal2 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER metal1 ;
  RECT 0.000 8.180 1.120 11.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 546.000 1076.880 549.540 1078.000 ;
  LAYER metal3 ;
  RECT 546.000 1076.880 549.540 1078.000 ;
  LAYER metal2 ;
  RECT 546.000 1076.880 549.540 1078.000 ;
  LAYER metal1 ;
  RECT 546.000 1076.880 549.540 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 537.320 1076.880 540.860 1078.000 ;
  LAYER metal3 ;
  RECT 537.320 1076.880 540.860 1078.000 ;
  LAYER metal2 ;
  RECT 537.320 1076.880 540.860 1078.000 ;
  LAYER metal1 ;
  RECT 537.320 1076.880 540.860 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 528.640 1076.880 532.180 1078.000 ;
  LAYER metal3 ;
  RECT 528.640 1076.880 532.180 1078.000 ;
  LAYER metal2 ;
  RECT 528.640 1076.880 532.180 1078.000 ;
  LAYER metal1 ;
  RECT 528.640 1076.880 532.180 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 485.240 1076.880 488.780 1078.000 ;
  LAYER metal3 ;
  RECT 485.240 1076.880 488.780 1078.000 ;
  LAYER metal2 ;
  RECT 485.240 1076.880 488.780 1078.000 ;
  LAYER metal1 ;
  RECT 485.240 1076.880 488.780 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 476.560 1076.880 480.100 1078.000 ;
  LAYER metal3 ;
  RECT 476.560 1076.880 480.100 1078.000 ;
  LAYER metal2 ;
  RECT 476.560 1076.880 480.100 1078.000 ;
  LAYER metal1 ;
  RECT 476.560 1076.880 480.100 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 467.880 1076.880 471.420 1078.000 ;
  LAYER metal3 ;
  RECT 467.880 1076.880 471.420 1078.000 ;
  LAYER metal2 ;
  RECT 467.880 1076.880 471.420 1078.000 ;
  LAYER metal1 ;
  RECT 467.880 1076.880 471.420 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 459.200 1076.880 462.740 1078.000 ;
  LAYER metal3 ;
  RECT 459.200 1076.880 462.740 1078.000 ;
  LAYER metal2 ;
  RECT 459.200 1076.880 462.740 1078.000 ;
  LAYER metal1 ;
  RECT 459.200 1076.880 462.740 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 450.520 1076.880 454.060 1078.000 ;
  LAYER metal3 ;
  RECT 450.520 1076.880 454.060 1078.000 ;
  LAYER metal2 ;
  RECT 450.520 1076.880 454.060 1078.000 ;
  LAYER metal1 ;
  RECT 450.520 1076.880 454.060 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 441.840 1076.880 445.380 1078.000 ;
  LAYER metal3 ;
  RECT 441.840 1076.880 445.380 1078.000 ;
  LAYER metal2 ;
  RECT 441.840 1076.880 445.380 1078.000 ;
  LAYER metal1 ;
  RECT 441.840 1076.880 445.380 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 398.440 1076.880 401.980 1078.000 ;
  LAYER metal3 ;
  RECT 398.440 1076.880 401.980 1078.000 ;
  LAYER metal2 ;
  RECT 398.440 1076.880 401.980 1078.000 ;
  LAYER metal1 ;
  RECT 398.440 1076.880 401.980 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 389.760 1076.880 393.300 1078.000 ;
  LAYER metal3 ;
  RECT 389.760 1076.880 393.300 1078.000 ;
  LAYER metal2 ;
  RECT 389.760 1076.880 393.300 1078.000 ;
  LAYER metal1 ;
  RECT 389.760 1076.880 393.300 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 381.080 1076.880 384.620 1078.000 ;
  LAYER metal3 ;
  RECT 381.080 1076.880 384.620 1078.000 ;
  LAYER metal2 ;
  RECT 381.080 1076.880 384.620 1078.000 ;
  LAYER metal1 ;
  RECT 381.080 1076.880 384.620 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 372.400 1076.880 375.940 1078.000 ;
  LAYER metal3 ;
  RECT 372.400 1076.880 375.940 1078.000 ;
  LAYER metal2 ;
  RECT 372.400 1076.880 375.940 1078.000 ;
  LAYER metal1 ;
  RECT 372.400 1076.880 375.940 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 363.720 1076.880 367.260 1078.000 ;
  LAYER metal3 ;
  RECT 363.720 1076.880 367.260 1078.000 ;
  LAYER metal2 ;
  RECT 363.720 1076.880 367.260 1078.000 ;
  LAYER metal1 ;
  RECT 363.720 1076.880 367.260 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 355.040 1076.880 358.580 1078.000 ;
  LAYER metal3 ;
  RECT 355.040 1076.880 358.580 1078.000 ;
  LAYER metal2 ;
  RECT 355.040 1076.880 358.580 1078.000 ;
  LAYER metal1 ;
  RECT 355.040 1076.880 358.580 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 311.640 1076.880 315.180 1078.000 ;
  LAYER metal3 ;
  RECT 311.640 1076.880 315.180 1078.000 ;
  LAYER metal2 ;
  RECT 311.640 1076.880 315.180 1078.000 ;
  LAYER metal1 ;
  RECT 311.640 1076.880 315.180 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 302.960 1076.880 306.500 1078.000 ;
  LAYER metal3 ;
  RECT 302.960 1076.880 306.500 1078.000 ;
  LAYER metal2 ;
  RECT 302.960 1076.880 306.500 1078.000 ;
  LAYER metal1 ;
  RECT 302.960 1076.880 306.500 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 294.280 1076.880 297.820 1078.000 ;
  LAYER metal3 ;
  RECT 294.280 1076.880 297.820 1078.000 ;
  LAYER metal2 ;
  RECT 294.280 1076.880 297.820 1078.000 ;
  LAYER metal1 ;
  RECT 294.280 1076.880 297.820 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 285.600 1076.880 289.140 1078.000 ;
  LAYER metal3 ;
  RECT 285.600 1076.880 289.140 1078.000 ;
  LAYER metal2 ;
  RECT 285.600 1076.880 289.140 1078.000 ;
  LAYER metal1 ;
  RECT 285.600 1076.880 289.140 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 276.920 1076.880 280.460 1078.000 ;
  LAYER metal3 ;
  RECT 276.920 1076.880 280.460 1078.000 ;
  LAYER metal2 ;
  RECT 276.920 1076.880 280.460 1078.000 ;
  LAYER metal1 ;
  RECT 276.920 1076.880 280.460 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 268.240 1076.880 271.780 1078.000 ;
  LAYER metal3 ;
  RECT 268.240 1076.880 271.780 1078.000 ;
  LAYER metal2 ;
  RECT 268.240 1076.880 271.780 1078.000 ;
  LAYER metal1 ;
  RECT 268.240 1076.880 271.780 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 224.840 1076.880 228.380 1078.000 ;
  LAYER metal3 ;
  RECT 224.840 1076.880 228.380 1078.000 ;
  LAYER metal2 ;
  RECT 224.840 1076.880 228.380 1078.000 ;
  LAYER metal1 ;
  RECT 224.840 1076.880 228.380 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 216.160 1076.880 219.700 1078.000 ;
  LAYER metal3 ;
  RECT 216.160 1076.880 219.700 1078.000 ;
  LAYER metal2 ;
  RECT 216.160 1076.880 219.700 1078.000 ;
  LAYER metal1 ;
  RECT 216.160 1076.880 219.700 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 207.480 1076.880 211.020 1078.000 ;
  LAYER metal3 ;
  RECT 207.480 1076.880 211.020 1078.000 ;
  LAYER metal2 ;
  RECT 207.480 1076.880 211.020 1078.000 ;
  LAYER metal1 ;
  RECT 207.480 1076.880 211.020 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 198.800 1076.880 202.340 1078.000 ;
  LAYER metal3 ;
  RECT 198.800 1076.880 202.340 1078.000 ;
  LAYER metal2 ;
  RECT 198.800 1076.880 202.340 1078.000 ;
  LAYER metal1 ;
  RECT 198.800 1076.880 202.340 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 190.120 1076.880 193.660 1078.000 ;
  LAYER metal3 ;
  RECT 190.120 1076.880 193.660 1078.000 ;
  LAYER metal2 ;
  RECT 190.120 1076.880 193.660 1078.000 ;
  LAYER metal1 ;
  RECT 190.120 1076.880 193.660 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 181.440 1076.880 184.980 1078.000 ;
  LAYER metal3 ;
  RECT 181.440 1076.880 184.980 1078.000 ;
  LAYER metal2 ;
  RECT 181.440 1076.880 184.980 1078.000 ;
  LAYER metal1 ;
  RECT 181.440 1076.880 184.980 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 138.040 1076.880 141.580 1078.000 ;
  LAYER metal3 ;
  RECT 138.040 1076.880 141.580 1078.000 ;
  LAYER metal2 ;
  RECT 138.040 1076.880 141.580 1078.000 ;
  LAYER metal1 ;
  RECT 138.040 1076.880 141.580 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 129.360 1076.880 132.900 1078.000 ;
  LAYER metal3 ;
  RECT 129.360 1076.880 132.900 1078.000 ;
  LAYER metal2 ;
  RECT 129.360 1076.880 132.900 1078.000 ;
  LAYER metal1 ;
  RECT 129.360 1076.880 132.900 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 120.680 1076.880 124.220 1078.000 ;
  LAYER metal3 ;
  RECT 120.680 1076.880 124.220 1078.000 ;
  LAYER metal2 ;
  RECT 120.680 1076.880 124.220 1078.000 ;
  LAYER metal1 ;
  RECT 120.680 1076.880 124.220 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 112.000 1076.880 115.540 1078.000 ;
  LAYER metal3 ;
  RECT 112.000 1076.880 115.540 1078.000 ;
  LAYER metal2 ;
  RECT 112.000 1076.880 115.540 1078.000 ;
  LAYER metal1 ;
  RECT 112.000 1076.880 115.540 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 103.320 1076.880 106.860 1078.000 ;
  LAYER metal3 ;
  RECT 103.320 1076.880 106.860 1078.000 ;
  LAYER metal2 ;
  RECT 103.320 1076.880 106.860 1078.000 ;
  LAYER metal1 ;
  RECT 103.320 1076.880 106.860 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 94.640 1076.880 98.180 1078.000 ;
  LAYER metal3 ;
  RECT 94.640 1076.880 98.180 1078.000 ;
  LAYER metal2 ;
  RECT 94.640 1076.880 98.180 1078.000 ;
  LAYER metal1 ;
  RECT 94.640 1076.880 98.180 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 51.240 1076.880 54.780 1078.000 ;
  LAYER metal3 ;
  RECT 51.240 1076.880 54.780 1078.000 ;
  LAYER metal2 ;
  RECT 51.240 1076.880 54.780 1078.000 ;
  LAYER metal1 ;
  RECT 51.240 1076.880 54.780 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 42.560 1076.880 46.100 1078.000 ;
  LAYER metal3 ;
  RECT 42.560 1076.880 46.100 1078.000 ;
  LAYER metal2 ;
  RECT 42.560 1076.880 46.100 1078.000 ;
  LAYER metal1 ;
  RECT 42.560 1076.880 46.100 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 33.880 1076.880 37.420 1078.000 ;
  LAYER metal3 ;
  RECT 33.880 1076.880 37.420 1078.000 ;
  LAYER metal2 ;
  RECT 33.880 1076.880 37.420 1078.000 ;
  LAYER metal1 ;
  RECT 33.880 1076.880 37.420 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 25.200 1076.880 28.740 1078.000 ;
  LAYER metal3 ;
  RECT 25.200 1076.880 28.740 1078.000 ;
  LAYER metal2 ;
  RECT 25.200 1076.880 28.740 1078.000 ;
  LAYER metal1 ;
  RECT 25.200 1076.880 28.740 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 16.520 1076.880 20.060 1078.000 ;
  LAYER metal3 ;
  RECT 16.520 1076.880 20.060 1078.000 ;
  LAYER metal2 ;
  RECT 16.520 1076.880 20.060 1078.000 ;
  LAYER metal1 ;
  RECT 16.520 1076.880 20.060 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 7.840 1076.880 11.380 1078.000 ;
  LAYER metal3 ;
  RECT 7.840 1076.880 11.380 1078.000 ;
  LAYER metal2 ;
  RECT 7.840 1076.880 11.380 1078.000 ;
  LAYER metal1 ;
  RECT 7.840 1076.880 11.380 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 543.520 0.000 547.060 1.120 ;
  LAYER metal3 ;
  RECT 543.520 0.000 547.060 1.120 ;
  LAYER metal2 ;
  RECT 543.520 0.000 547.060 1.120 ;
  LAYER metal1 ;
  RECT 543.520 0.000 547.060 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 522.440 0.000 525.980 1.120 ;
  LAYER metal3 ;
  RECT 522.440 0.000 525.980 1.120 ;
  LAYER metal2 ;
  RECT 522.440 0.000 525.980 1.120 ;
  LAYER metal1 ;
  RECT 522.440 0.000 525.980 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 500.740 0.000 504.280 1.120 ;
  LAYER metal3 ;
  RECT 500.740 0.000 504.280 1.120 ;
  LAYER metal2 ;
  RECT 500.740 0.000 504.280 1.120 ;
  LAYER metal1 ;
  RECT 500.740 0.000 504.280 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 474.080 0.000 477.620 1.120 ;
  LAYER metal3 ;
  RECT 474.080 0.000 477.620 1.120 ;
  LAYER metal2 ;
  RECT 474.080 0.000 477.620 1.120 ;
  LAYER metal1 ;
  RECT 474.080 0.000 477.620 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 457.340 0.000 460.880 1.120 ;
  LAYER metal3 ;
  RECT 457.340 0.000 460.880 1.120 ;
  LAYER metal2 ;
  RECT 457.340 0.000 460.880 1.120 ;
  LAYER metal1 ;
  RECT 457.340 0.000 460.880 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 344.500 0.000 348.040 1.120 ;
  LAYER metal3 ;
  RECT 344.500 0.000 348.040 1.120 ;
  LAYER metal2 ;
  RECT 344.500 0.000 348.040 1.120 ;
  LAYER metal1 ;
  RECT 344.500 0.000 348.040 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 308.540 0.000 312.080 1.120 ;
  LAYER metal3 ;
  RECT 308.540 0.000 312.080 1.120 ;
  LAYER metal2 ;
  RECT 308.540 0.000 312.080 1.120 ;
  LAYER metal1 ;
  RECT 308.540 0.000 312.080 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 299.860 0.000 303.400 1.120 ;
  LAYER metal3 ;
  RECT 299.860 0.000 303.400 1.120 ;
  LAYER metal2 ;
  RECT 299.860 0.000 303.400 1.120 ;
  LAYER metal1 ;
  RECT 299.860 0.000 303.400 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 278.160 0.000 281.700 1.120 ;
  LAYER metal3 ;
  RECT 278.160 0.000 281.700 1.120 ;
  LAYER metal2 ;
  RECT 278.160 0.000 281.700 1.120 ;
  LAYER metal1 ;
  RECT 278.160 0.000 281.700 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 257.080 0.000 260.620 1.120 ;
  LAYER metal3 ;
  RECT 257.080 0.000 260.620 1.120 ;
  LAYER metal2 ;
  RECT 257.080 0.000 260.620 1.120 ;
  LAYER metal1 ;
  RECT 257.080 0.000 260.620 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 235.380 0.000 238.920 1.120 ;
  LAYER metal3 ;
  RECT 235.380 0.000 238.920 1.120 ;
  LAYER metal2 ;
  RECT 235.380 0.000 238.920 1.120 ;
  LAYER metal1 ;
  RECT 235.380 0.000 238.920 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER metal3 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER metal2 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER metal1 ;
  RECT 126.880 0.000 130.420 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER metal3 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER metal2 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER metal1 ;
  RECT 100.220 0.000 103.760 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER metal3 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER metal2 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER metal1 ;
  RECT 83.480 0.000 87.020 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER metal3 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER metal2 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER metal1 ;
  RECT 56.820 0.000 60.360 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal3 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal2 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER metal1 ;
  RECT 35.740 0.000 39.280 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER metal3 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER metal2 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER metal1 ;
  RECT 14.040 0.000 17.580 1.120 ;
 END
END VCC
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER metal4 ;
  RECT 562.460 1062.660 563.580 1065.900 ;
  LAYER metal3 ;
  RECT 562.460 1062.660 563.580 1065.900 ;
  LAYER metal2 ;
  RECT 562.460 1062.660 563.580 1065.900 ;
  LAYER metal1 ;
  RECT 562.460 1062.660 563.580 1065.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 1054.820 563.580 1058.060 ;
  LAYER metal3 ;
  RECT 562.460 1054.820 563.580 1058.060 ;
  LAYER metal2 ;
  RECT 562.460 1054.820 563.580 1058.060 ;
  LAYER metal1 ;
  RECT 562.460 1054.820 563.580 1058.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 1046.980 563.580 1050.220 ;
  LAYER metal3 ;
  RECT 562.460 1046.980 563.580 1050.220 ;
  LAYER metal2 ;
  RECT 562.460 1046.980 563.580 1050.220 ;
  LAYER metal1 ;
  RECT 562.460 1046.980 563.580 1050.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 1039.140 563.580 1042.380 ;
  LAYER metal3 ;
  RECT 562.460 1039.140 563.580 1042.380 ;
  LAYER metal2 ;
  RECT 562.460 1039.140 563.580 1042.380 ;
  LAYER metal1 ;
  RECT 562.460 1039.140 563.580 1042.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 1031.300 563.580 1034.540 ;
  LAYER metal3 ;
  RECT 562.460 1031.300 563.580 1034.540 ;
  LAYER metal2 ;
  RECT 562.460 1031.300 563.580 1034.540 ;
  LAYER metal1 ;
  RECT 562.460 1031.300 563.580 1034.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 992.100 563.580 995.340 ;
  LAYER metal3 ;
  RECT 562.460 992.100 563.580 995.340 ;
  LAYER metal2 ;
  RECT 562.460 992.100 563.580 995.340 ;
  LAYER metal1 ;
  RECT 562.460 992.100 563.580 995.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 984.260 563.580 987.500 ;
  LAYER metal3 ;
  RECT 562.460 984.260 563.580 987.500 ;
  LAYER metal2 ;
  RECT 562.460 984.260 563.580 987.500 ;
  LAYER metal1 ;
  RECT 562.460 984.260 563.580 987.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 976.420 563.580 979.660 ;
  LAYER metal3 ;
  RECT 562.460 976.420 563.580 979.660 ;
  LAYER metal2 ;
  RECT 562.460 976.420 563.580 979.660 ;
  LAYER metal1 ;
  RECT 562.460 976.420 563.580 979.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 968.580 563.580 971.820 ;
  LAYER metal3 ;
  RECT 562.460 968.580 563.580 971.820 ;
  LAYER metal2 ;
  RECT 562.460 968.580 563.580 971.820 ;
  LAYER metal1 ;
  RECT 562.460 968.580 563.580 971.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 960.740 563.580 963.980 ;
  LAYER metal3 ;
  RECT 562.460 960.740 563.580 963.980 ;
  LAYER metal2 ;
  RECT 562.460 960.740 563.580 963.980 ;
  LAYER metal1 ;
  RECT 562.460 960.740 563.580 963.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 952.900 563.580 956.140 ;
  LAYER metal3 ;
  RECT 562.460 952.900 563.580 956.140 ;
  LAYER metal2 ;
  RECT 562.460 952.900 563.580 956.140 ;
  LAYER metal1 ;
  RECT 562.460 952.900 563.580 956.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 913.700 563.580 916.940 ;
  LAYER metal3 ;
  RECT 562.460 913.700 563.580 916.940 ;
  LAYER metal2 ;
  RECT 562.460 913.700 563.580 916.940 ;
  LAYER metal1 ;
  RECT 562.460 913.700 563.580 916.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 905.860 563.580 909.100 ;
  LAYER metal3 ;
  RECT 562.460 905.860 563.580 909.100 ;
  LAYER metal2 ;
  RECT 562.460 905.860 563.580 909.100 ;
  LAYER metal1 ;
  RECT 562.460 905.860 563.580 909.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 898.020 563.580 901.260 ;
  LAYER metal3 ;
  RECT 562.460 898.020 563.580 901.260 ;
  LAYER metal2 ;
  RECT 562.460 898.020 563.580 901.260 ;
  LAYER metal1 ;
  RECT 562.460 898.020 563.580 901.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 890.180 563.580 893.420 ;
  LAYER metal3 ;
  RECT 562.460 890.180 563.580 893.420 ;
  LAYER metal2 ;
  RECT 562.460 890.180 563.580 893.420 ;
  LAYER metal1 ;
  RECT 562.460 890.180 563.580 893.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 882.340 563.580 885.580 ;
  LAYER metal3 ;
  RECT 562.460 882.340 563.580 885.580 ;
  LAYER metal2 ;
  RECT 562.460 882.340 563.580 885.580 ;
  LAYER metal1 ;
  RECT 562.460 882.340 563.580 885.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 874.500 563.580 877.740 ;
  LAYER metal3 ;
  RECT 562.460 874.500 563.580 877.740 ;
  LAYER metal2 ;
  RECT 562.460 874.500 563.580 877.740 ;
  LAYER metal1 ;
  RECT 562.460 874.500 563.580 877.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 835.300 563.580 838.540 ;
  LAYER metal3 ;
  RECT 562.460 835.300 563.580 838.540 ;
  LAYER metal2 ;
  RECT 562.460 835.300 563.580 838.540 ;
  LAYER metal1 ;
  RECT 562.460 835.300 563.580 838.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 827.460 563.580 830.700 ;
  LAYER metal3 ;
  RECT 562.460 827.460 563.580 830.700 ;
  LAYER metal2 ;
  RECT 562.460 827.460 563.580 830.700 ;
  LAYER metal1 ;
  RECT 562.460 827.460 563.580 830.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 819.620 563.580 822.860 ;
  LAYER metal3 ;
  RECT 562.460 819.620 563.580 822.860 ;
  LAYER metal2 ;
  RECT 562.460 819.620 563.580 822.860 ;
  LAYER metal1 ;
  RECT 562.460 819.620 563.580 822.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 811.780 563.580 815.020 ;
  LAYER metal3 ;
  RECT 562.460 811.780 563.580 815.020 ;
  LAYER metal2 ;
  RECT 562.460 811.780 563.580 815.020 ;
  LAYER metal1 ;
  RECT 562.460 811.780 563.580 815.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 803.940 563.580 807.180 ;
  LAYER metal3 ;
  RECT 562.460 803.940 563.580 807.180 ;
  LAYER metal2 ;
  RECT 562.460 803.940 563.580 807.180 ;
  LAYER metal1 ;
  RECT 562.460 803.940 563.580 807.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 796.100 563.580 799.340 ;
  LAYER metal3 ;
  RECT 562.460 796.100 563.580 799.340 ;
  LAYER metal2 ;
  RECT 562.460 796.100 563.580 799.340 ;
  LAYER metal1 ;
  RECT 562.460 796.100 563.580 799.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 756.900 563.580 760.140 ;
  LAYER metal3 ;
  RECT 562.460 756.900 563.580 760.140 ;
  LAYER metal2 ;
  RECT 562.460 756.900 563.580 760.140 ;
  LAYER metal1 ;
  RECT 562.460 756.900 563.580 760.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 749.060 563.580 752.300 ;
  LAYER metal3 ;
  RECT 562.460 749.060 563.580 752.300 ;
  LAYER metal2 ;
  RECT 562.460 749.060 563.580 752.300 ;
  LAYER metal1 ;
  RECT 562.460 749.060 563.580 752.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 741.220 563.580 744.460 ;
  LAYER metal3 ;
  RECT 562.460 741.220 563.580 744.460 ;
  LAYER metal2 ;
  RECT 562.460 741.220 563.580 744.460 ;
  LAYER metal1 ;
  RECT 562.460 741.220 563.580 744.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 733.380 563.580 736.620 ;
  LAYER metal3 ;
  RECT 562.460 733.380 563.580 736.620 ;
  LAYER metal2 ;
  RECT 562.460 733.380 563.580 736.620 ;
  LAYER metal1 ;
  RECT 562.460 733.380 563.580 736.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 725.540 563.580 728.780 ;
  LAYER metal3 ;
  RECT 562.460 725.540 563.580 728.780 ;
  LAYER metal2 ;
  RECT 562.460 725.540 563.580 728.780 ;
  LAYER metal1 ;
  RECT 562.460 725.540 563.580 728.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 717.700 563.580 720.940 ;
  LAYER metal3 ;
  RECT 562.460 717.700 563.580 720.940 ;
  LAYER metal2 ;
  RECT 562.460 717.700 563.580 720.940 ;
  LAYER metal1 ;
  RECT 562.460 717.700 563.580 720.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 678.500 563.580 681.740 ;
  LAYER metal3 ;
  RECT 562.460 678.500 563.580 681.740 ;
  LAYER metal2 ;
  RECT 562.460 678.500 563.580 681.740 ;
  LAYER metal1 ;
  RECT 562.460 678.500 563.580 681.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 670.660 563.580 673.900 ;
  LAYER metal3 ;
  RECT 562.460 670.660 563.580 673.900 ;
  LAYER metal2 ;
  RECT 562.460 670.660 563.580 673.900 ;
  LAYER metal1 ;
  RECT 562.460 670.660 563.580 673.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 662.820 563.580 666.060 ;
  LAYER metal3 ;
  RECT 562.460 662.820 563.580 666.060 ;
  LAYER metal2 ;
  RECT 562.460 662.820 563.580 666.060 ;
  LAYER metal1 ;
  RECT 562.460 662.820 563.580 666.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 654.980 563.580 658.220 ;
  LAYER metal3 ;
  RECT 562.460 654.980 563.580 658.220 ;
  LAYER metal2 ;
  RECT 562.460 654.980 563.580 658.220 ;
  LAYER metal1 ;
  RECT 562.460 654.980 563.580 658.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 647.140 563.580 650.380 ;
  LAYER metal3 ;
  RECT 562.460 647.140 563.580 650.380 ;
  LAYER metal2 ;
  RECT 562.460 647.140 563.580 650.380 ;
  LAYER metal1 ;
  RECT 562.460 647.140 563.580 650.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 639.300 563.580 642.540 ;
  LAYER metal3 ;
  RECT 562.460 639.300 563.580 642.540 ;
  LAYER metal2 ;
  RECT 562.460 639.300 563.580 642.540 ;
  LAYER metal1 ;
  RECT 562.460 639.300 563.580 642.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 600.100 563.580 603.340 ;
  LAYER metal3 ;
  RECT 562.460 600.100 563.580 603.340 ;
  LAYER metal2 ;
  RECT 562.460 600.100 563.580 603.340 ;
  LAYER metal1 ;
  RECT 562.460 600.100 563.580 603.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 592.260 563.580 595.500 ;
  LAYER metal3 ;
  RECT 562.460 592.260 563.580 595.500 ;
  LAYER metal2 ;
  RECT 562.460 592.260 563.580 595.500 ;
  LAYER metal1 ;
  RECT 562.460 592.260 563.580 595.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 584.420 563.580 587.660 ;
  LAYER metal3 ;
  RECT 562.460 584.420 563.580 587.660 ;
  LAYER metal2 ;
  RECT 562.460 584.420 563.580 587.660 ;
  LAYER metal1 ;
  RECT 562.460 584.420 563.580 587.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 576.580 563.580 579.820 ;
  LAYER metal3 ;
  RECT 562.460 576.580 563.580 579.820 ;
  LAYER metal2 ;
  RECT 562.460 576.580 563.580 579.820 ;
  LAYER metal1 ;
  RECT 562.460 576.580 563.580 579.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 568.740 563.580 571.980 ;
  LAYER metal3 ;
  RECT 562.460 568.740 563.580 571.980 ;
  LAYER metal2 ;
  RECT 562.460 568.740 563.580 571.980 ;
  LAYER metal1 ;
  RECT 562.460 568.740 563.580 571.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 560.900 563.580 564.140 ;
  LAYER metal3 ;
  RECT 562.460 560.900 563.580 564.140 ;
  LAYER metal2 ;
  RECT 562.460 560.900 563.580 564.140 ;
  LAYER metal1 ;
  RECT 562.460 560.900 563.580 564.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 521.700 563.580 524.940 ;
  LAYER metal3 ;
  RECT 562.460 521.700 563.580 524.940 ;
  LAYER metal2 ;
  RECT 562.460 521.700 563.580 524.940 ;
  LAYER metal1 ;
  RECT 562.460 521.700 563.580 524.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 513.860 563.580 517.100 ;
  LAYER metal3 ;
  RECT 562.460 513.860 563.580 517.100 ;
  LAYER metal2 ;
  RECT 562.460 513.860 563.580 517.100 ;
  LAYER metal1 ;
  RECT 562.460 513.860 563.580 517.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 506.020 563.580 509.260 ;
  LAYER metal3 ;
  RECT 562.460 506.020 563.580 509.260 ;
  LAYER metal2 ;
  RECT 562.460 506.020 563.580 509.260 ;
  LAYER metal1 ;
  RECT 562.460 506.020 563.580 509.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 498.180 563.580 501.420 ;
  LAYER metal3 ;
  RECT 562.460 498.180 563.580 501.420 ;
  LAYER metal2 ;
  RECT 562.460 498.180 563.580 501.420 ;
  LAYER metal1 ;
  RECT 562.460 498.180 563.580 501.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 490.340 563.580 493.580 ;
  LAYER metal3 ;
  RECT 562.460 490.340 563.580 493.580 ;
  LAYER metal2 ;
  RECT 562.460 490.340 563.580 493.580 ;
  LAYER metal1 ;
  RECT 562.460 490.340 563.580 493.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 482.500 563.580 485.740 ;
  LAYER metal3 ;
  RECT 562.460 482.500 563.580 485.740 ;
  LAYER metal2 ;
  RECT 562.460 482.500 563.580 485.740 ;
  LAYER metal1 ;
  RECT 562.460 482.500 563.580 485.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 443.300 563.580 446.540 ;
  LAYER metal3 ;
  RECT 562.460 443.300 563.580 446.540 ;
  LAYER metal2 ;
  RECT 562.460 443.300 563.580 446.540 ;
  LAYER metal1 ;
  RECT 562.460 443.300 563.580 446.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 435.460 563.580 438.700 ;
  LAYER metal3 ;
  RECT 562.460 435.460 563.580 438.700 ;
  LAYER metal2 ;
  RECT 562.460 435.460 563.580 438.700 ;
  LAYER metal1 ;
  RECT 562.460 435.460 563.580 438.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 427.620 563.580 430.860 ;
  LAYER metal3 ;
  RECT 562.460 427.620 563.580 430.860 ;
  LAYER metal2 ;
  RECT 562.460 427.620 563.580 430.860 ;
  LAYER metal1 ;
  RECT 562.460 427.620 563.580 430.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 419.780 563.580 423.020 ;
  LAYER metal3 ;
  RECT 562.460 419.780 563.580 423.020 ;
  LAYER metal2 ;
  RECT 562.460 419.780 563.580 423.020 ;
  LAYER metal1 ;
  RECT 562.460 419.780 563.580 423.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 411.940 563.580 415.180 ;
  LAYER metal3 ;
  RECT 562.460 411.940 563.580 415.180 ;
  LAYER metal2 ;
  RECT 562.460 411.940 563.580 415.180 ;
  LAYER metal1 ;
  RECT 562.460 411.940 563.580 415.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 404.100 563.580 407.340 ;
  LAYER metal3 ;
  RECT 562.460 404.100 563.580 407.340 ;
  LAYER metal2 ;
  RECT 562.460 404.100 563.580 407.340 ;
  LAYER metal1 ;
  RECT 562.460 404.100 563.580 407.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 364.900 563.580 368.140 ;
  LAYER metal3 ;
  RECT 562.460 364.900 563.580 368.140 ;
  LAYER metal2 ;
  RECT 562.460 364.900 563.580 368.140 ;
  LAYER metal1 ;
  RECT 562.460 364.900 563.580 368.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 357.060 563.580 360.300 ;
  LAYER metal3 ;
  RECT 562.460 357.060 563.580 360.300 ;
  LAYER metal2 ;
  RECT 562.460 357.060 563.580 360.300 ;
  LAYER metal1 ;
  RECT 562.460 357.060 563.580 360.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 349.220 563.580 352.460 ;
  LAYER metal3 ;
  RECT 562.460 349.220 563.580 352.460 ;
  LAYER metal2 ;
  RECT 562.460 349.220 563.580 352.460 ;
  LAYER metal1 ;
  RECT 562.460 349.220 563.580 352.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 341.380 563.580 344.620 ;
  LAYER metal3 ;
  RECT 562.460 341.380 563.580 344.620 ;
  LAYER metal2 ;
  RECT 562.460 341.380 563.580 344.620 ;
  LAYER metal1 ;
  RECT 562.460 341.380 563.580 344.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 333.540 563.580 336.780 ;
  LAYER metal3 ;
  RECT 562.460 333.540 563.580 336.780 ;
  LAYER metal2 ;
  RECT 562.460 333.540 563.580 336.780 ;
  LAYER metal1 ;
  RECT 562.460 333.540 563.580 336.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 325.700 563.580 328.940 ;
  LAYER metal3 ;
  RECT 562.460 325.700 563.580 328.940 ;
  LAYER metal2 ;
  RECT 562.460 325.700 563.580 328.940 ;
  LAYER metal1 ;
  RECT 562.460 325.700 563.580 328.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 286.500 563.580 289.740 ;
  LAYER metal3 ;
  RECT 562.460 286.500 563.580 289.740 ;
  LAYER metal2 ;
  RECT 562.460 286.500 563.580 289.740 ;
  LAYER metal1 ;
  RECT 562.460 286.500 563.580 289.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 278.660 563.580 281.900 ;
  LAYER metal3 ;
  RECT 562.460 278.660 563.580 281.900 ;
  LAYER metal2 ;
  RECT 562.460 278.660 563.580 281.900 ;
  LAYER metal1 ;
  RECT 562.460 278.660 563.580 281.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 270.820 563.580 274.060 ;
  LAYER metal3 ;
  RECT 562.460 270.820 563.580 274.060 ;
  LAYER metal2 ;
  RECT 562.460 270.820 563.580 274.060 ;
  LAYER metal1 ;
  RECT 562.460 270.820 563.580 274.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 262.980 563.580 266.220 ;
  LAYER metal3 ;
  RECT 562.460 262.980 563.580 266.220 ;
  LAYER metal2 ;
  RECT 562.460 262.980 563.580 266.220 ;
  LAYER metal1 ;
  RECT 562.460 262.980 563.580 266.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 255.140 563.580 258.380 ;
  LAYER metal3 ;
  RECT 562.460 255.140 563.580 258.380 ;
  LAYER metal2 ;
  RECT 562.460 255.140 563.580 258.380 ;
  LAYER metal1 ;
  RECT 562.460 255.140 563.580 258.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 247.300 563.580 250.540 ;
  LAYER metal3 ;
  RECT 562.460 247.300 563.580 250.540 ;
  LAYER metal2 ;
  RECT 562.460 247.300 563.580 250.540 ;
  LAYER metal1 ;
  RECT 562.460 247.300 563.580 250.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 208.100 563.580 211.340 ;
  LAYER metal3 ;
  RECT 562.460 208.100 563.580 211.340 ;
  LAYER metal2 ;
  RECT 562.460 208.100 563.580 211.340 ;
  LAYER metal1 ;
  RECT 562.460 208.100 563.580 211.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 200.260 563.580 203.500 ;
  LAYER metal3 ;
  RECT 562.460 200.260 563.580 203.500 ;
  LAYER metal2 ;
  RECT 562.460 200.260 563.580 203.500 ;
  LAYER metal1 ;
  RECT 562.460 200.260 563.580 203.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 192.420 563.580 195.660 ;
  LAYER metal3 ;
  RECT 562.460 192.420 563.580 195.660 ;
  LAYER metal2 ;
  RECT 562.460 192.420 563.580 195.660 ;
  LAYER metal1 ;
  RECT 562.460 192.420 563.580 195.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 184.580 563.580 187.820 ;
  LAYER metal3 ;
  RECT 562.460 184.580 563.580 187.820 ;
  LAYER metal2 ;
  RECT 562.460 184.580 563.580 187.820 ;
  LAYER metal1 ;
  RECT 562.460 184.580 563.580 187.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 176.740 563.580 179.980 ;
  LAYER metal3 ;
  RECT 562.460 176.740 563.580 179.980 ;
  LAYER metal2 ;
  RECT 562.460 176.740 563.580 179.980 ;
  LAYER metal1 ;
  RECT 562.460 176.740 563.580 179.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 168.900 563.580 172.140 ;
  LAYER metal3 ;
  RECT 562.460 168.900 563.580 172.140 ;
  LAYER metal2 ;
  RECT 562.460 168.900 563.580 172.140 ;
  LAYER metal1 ;
  RECT 562.460 168.900 563.580 172.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 129.700 563.580 132.940 ;
  LAYER metal3 ;
  RECT 562.460 129.700 563.580 132.940 ;
  LAYER metal2 ;
  RECT 562.460 129.700 563.580 132.940 ;
  LAYER metal1 ;
  RECT 562.460 129.700 563.580 132.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 121.860 563.580 125.100 ;
  LAYER metal3 ;
  RECT 562.460 121.860 563.580 125.100 ;
  LAYER metal2 ;
  RECT 562.460 121.860 563.580 125.100 ;
  LAYER metal1 ;
  RECT 562.460 121.860 563.580 125.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 114.020 563.580 117.260 ;
  LAYER metal3 ;
  RECT 562.460 114.020 563.580 117.260 ;
  LAYER metal2 ;
  RECT 562.460 114.020 563.580 117.260 ;
  LAYER metal1 ;
  RECT 562.460 114.020 563.580 117.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 106.180 563.580 109.420 ;
  LAYER metal3 ;
  RECT 562.460 106.180 563.580 109.420 ;
  LAYER metal2 ;
  RECT 562.460 106.180 563.580 109.420 ;
  LAYER metal1 ;
  RECT 562.460 106.180 563.580 109.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 98.340 563.580 101.580 ;
  LAYER metal3 ;
  RECT 562.460 98.340 563.580 101.580 ;
  LAYER metal2 ;
  RECT 562.460 98.340 563.580 101.580 ;
  LAYER metal1 ;
  RECT 562.460 98.340 563.580 101.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 90.500 563.580 93.740 ;
  LAYER metal3 ;
  RECT 562.460 90.500 563.580 93.740 ;
  LAYER metal2 ;
  RECT 562.460 90.500 563.580 93.740 ;
  LAYER metal1 ;
  RECT 562.460 90.500 563.580 93.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 51.300 563.580 54.540 ;
  LAYER metal3 ;
  RECT 562.460 51.300 563.580 54.540 ;
  LAYER metal2 ;
  RECT 562.460 51.300 563.580 54.540 ;
  LAYER metal1 ;
  RECT 562.460 51.300 563.580 54.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 43.460 563.580 46.700 ;
  LAYER metal3 ;
  RECT 562.460 43.460 563.580 46.700 ;
  LAYER metal2 ;
  RECT 562.460 43.460 563.580 46.700 ;
  LAYER metal1 ;
  RECT 562.460 43.460 563.580 46.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 35.620 563.580 38.860 ;
  LAYER metal3 ;
  RECT 562.460 35.620 563.580 38.860 ;
  LAYER metal2 ;
  RECT 562.460 35.620 563.580 38.860 ;
  LAYER metal1 ;
  RECT 562.460 35.620 563.580 38.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 27.780 563.580 31.020 ;
  LAYER metal3 ;
  RECT 562.460 27.780 563.580 31.020 ;
  LAYER metal2 ;
  RECT 562.460 27.780 563.580 31.020 ;
  LAYER metal1 ;
  RECT 562.460 27.780 563.580 31.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 19.940 563.580 23.180 ;
  LAYER metal3 ;
  RECT 562.460 19.940 563.580 23.180 ;
  LAYER metal2 ;
  RECT 562.460 19.940 563.580 23.180 ;
  LAYER metal1 ;
  RECT 562.460 19.940 563.580 23.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 562.460 12.100 563.580 15.340 ;
  LAYER metal3 ;
  RECT 562.460 12.100 563.580 15.340 ;
  LAYER metal2 ;
  RECT 562.460 12.100 563.580 15.340 ;
  LAYER metal1 ;
  RECT 562.460 12.100 563.580 15.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1062.660 1.120 1065.900 ;
  LAYER metal3 ;
  RECT 0.000 1062.660 1.120 1065.900 ;
  LAYER metal2 ;
  RECT 0.000 1062.660 1.120 1065.900 ;
  LAYER metal1 ;
  RECT 0.000 1062.660 1.120 1065.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1054.820 1.120 1058.060 ;
  LAYER metal3 ;
  RECT 0.000 1054.820 1.120 1058.060 ;
  LAYER metal2 ;
  RECT 0.000 1054.820 1.120 1058.060 ;
  LAYER metal1 ;
  RECT 0.000 1054.820 1.120 1058.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1046.980 1.120 1050.220 ;
  LAYER metal3 ;
  RECT 0.000 1046.980 1.120 1050.220 ;
  LAYER metal2 ;
  RECT 0.000 1046.980 1.120 1050.220 ;
  LAYER metal1 ;
  RECT 0.000 1046.980 1.120 1050.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1039.140 1.120 1042.380 ;
  LAYER metal3 ;
  RECT 0.000 1039.140 1.120 1042.380 ;
  LAYER metal2 ;
  RECT 0.000 1039.140 1.120 1042.380 ;
  LAYER metal1 ;
  RECT 0.000 1039.140 1.120 1042.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 1031.300 1.120 1034.540 ;
  LAYER metal3 ;
  RECT 0.000 1031.300 1.120 1034.540 ;
  LAYER metal2 ;
  RECT 0.000 1031.300 1.120 1034.540 ;
  LAYER metal1 ;
  RECT 0.000 1031.300 1.120 1034.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 992.100 1.120 995.340 ;
  LAYER metal3 ;
  RECT 0.000 992.100 1.120 995.340 ;
  LAYER metal2 ;
  RECT 0.000 992.100 1.120 995.340 ;
  LAYER metal1 ;
  RECT 0.000 992.100 1.120 995.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 984.260 1.120 987.500 ;
  LAYER metal3 ;
  RECT 0.000 984.260 1.120 987.500 ;
  LAYER metal2 ;
  RECT 0.000 984.260 1.120 987.500 ;
  LAYER metal1 ;
  RECT 0.000 984.260 1.120 987.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 976.420 1.120 979.660 ;
  LAYER metal3 ;
  RECT 0.000 976.420 1.120 979.660 ;
  LAYER metal2 ;
  RECT 0.000 976.420 1.120 979.660 ;
  LAYER metal1 ;
  RECT 0.000 976.420 1.120 979.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 968.580 1.120 971.820 ;
  LAYER metal3 ;
  RECT 0.000 968.580 1.120 971.820 ;
  LAYER metal2 ;
  RECT 0.000 968.580 1.120 971.820 ;
  LAYER metal1 ;
  RECT 0.000 968.580 1.120 971.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 960.740 1.120 963.980 ;
  LAYER metal3 ;
  RECT 0.000 960.740 1.120 963.980 ;
  LAYER metal2 ;
  RECT 0.000 960.740 1.120 963.980 ;
  LAYER metal1 ;
  RECT 0.000 960.740 1.120 963.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 952.900 1.120 956.140 ;
  LAYER metal3 ;
  RECT 0.000 952.900 1.120 956.140 ;
  LAYER metal2 ;
  RECT 0.000 952.900 1.120 956.140 ;
  LAYER metal1 ;
  RECT 0.000 952.900 1.120 956.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 913.700 1.120 916.940 ;
  LAYER metal3 ;
  RECT 0.000 913.700 1.120 916.940 ;
  LAYER metal2 ;
  RECT 0.000 913.700 1.120 916.940 ;
  LAYER metal1 ;
  RECT 0.000 913.700 1.120 916.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 905.860 1.120 909.100 ;
  LAYER metal3 ;
  RECT 0.000 905.860 1.120 909.100 ;
  LAYER metal2 ;
  RECT 0.000 905.860 1.120 909.100 ;
  LAYER metal1 ;
  RECT 0.000 905.860 1.120 909.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 898.020 1.120 901.260 ;
  LAYER metal3 ;
  RECT 0.000 898.020 1.120 901.260 ;
  LAYER metal2 ;
  RECT 0.000 898.020 1.120 901.260 ;
  LAYER metal1 ;
  RECT 0.000 898.020 1.120 901.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 890.180 1.120 893.420 ;
  LAYER metal3 ;
  RECT 0.000 890.180 1.120 893.420 ;
  LAYER metal2 ;
  RECT 0.000 890.180 1.120 893.420 ;
  LAYER metal1 ;
  RECT 0.000 890.180 1.120 893.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 882.340 1.120 885.580 ;
  LAYER metal3 ;
  RECT 0.000 882.340 1.120 885.580 ;
  LAYER metal2 ;
  RECT 0.000 882.340 1.120 885.580 ;
  LAYER metal1 ;
  RECT 0.000 882.340 1.120 885.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 874.500 1.120 877.740 ;
  LAYER metal3 ;
  RECT 0.000 874.500 1.120 877.740 ;
  LAYER metal2 ;
  RECT 0.000 874.500 1.120 877.740 ;
  LAYER metal1 ;
  RECT 0.000 874.500 1.120 877.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 835.300 1.120 838.540 ;
  LAYER metal3 ;
  RECT 0.000 835.300 1.120 838.540 ;
  LAYER metal2 ;
  RECT 0.000 835.300 1.120 838.540 ;
  LAYER metal1 ;
  RECT 0.000 835.300 1.120 838.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 827.460 1.120 830.700 ;
  LAYER metal3 ;
  RECT 0.000 827.460 1.120 830.700 ;
  LAYER metal2 ;
  RECT 0.000 827.460 1.120 830.700 ;
  LAYER metal1 ;
  RECT 0.000 827.460 1.120 830.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 819.620 1.120 822.860 ;
  LAYER metal3 ;
  RECT 0.000 819.620 1.120 822.860 ;
  LAYER metal2 ;
  RECT 0.000 819.620 1.120 822.860 ;
  LAYER metal1 ;
  RECT 0.000 819.620 1.120 822.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 811.780 1.120 815.020 ;
  LAYER metal3 ;
  RECT 0.000 811.780 1.120 815.020 ;
  LAYER metal2 ;
  RECT 0.000 811.780 1.120 815.020 ;
  LAYER metal1 ;
  RECT 0.000 811.780 1.120 815.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 803.940 1.120 807.180 ;
  LAYER metal3 ;
  RECT 0.000 803.940 1.120 807.180 ;
  LAYER metal2 ;
  RECT 0.000 803.940 1.120 807.180 ;
  LAYER metal1 ;
  RECT 0.000 803.940 1.120 807.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 796.100 1.120 799.340 ;
  LAYER metal3 ;
  RECT 0.000 796.100 1.120 799.340 ;
  LAYER metal2 ;
  RECT 0.000 796.100 1.120 799.340 ;
  LAYER metal1 ;
  RECT 0.000 796.100 1.120 799.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 756.900 1.120 760.140 ;
  LAYER metal3 ;
  RECT 0.000 756.900 1.120 760.140 ;
  LAYER metal2 ;
  RECT 0.000 756.900 1.120 760.140 ;
  LAYER metal1 ;
  RECT 0.000 756.900 1.120 760.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 749.060 1.120 752.300 ;
  LAYER metal3 ;
  RECT 0.000 749.060 1.120 752.300 ;
  LAYER metal2 ;
  RECT 0.000 749.060 1.120 752.300 ;
  LAYER metal1 ;
  RECT 0.000 749.060 1.120 752.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 741.220 1.120 744.460 ;
  LAYER metal3 ;
  RECT 0.000 741.220 1.120 744.460 ;
  LAYER metal2 ;
  RECT 0.000 741.220 1.120 744.460 ;
  LAYER metal1 ;
  RECT 0.000 741.220 1.120 744.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 733.380 1.120 736.620 ;
  LAYER metal3 ;
  RECT 0.000 733.380 1.120 736.620 ;
  LAYER metal2 ;
  RECT 0.000 733.380 1.120 736.620 ;
  LAYER metal1 ;
  RECT 0.000 733.380 1.120 736.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 725.540 1.120 728.780 ;
  LAYER metal3 ;
  RECT 0.000 725.540 1.120 728.780 ;
  LAYER metal2 ;
  RECT 0.000 725.540 1.120 728.780 ;
  LAYER metal1 ;
  RECT 0.000 725.540 1.120 728.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 717.700 1.120 720.940 ;
  LAYER metal3 ;
  RECT 0.000 717.700 1.120 720.940 ;
  LAYER metal2 ;
  RECT 0.000 717.700 1.120 720.940 ;
  LAYER metal1 ;
  RECT 0.000 717.700 1.120 720.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 678.500 1.120 681.740 ;
  LAYER metal3 ;
  RECT 0.000 678.500 1.120 681.740 ;
  LAYER metal2 ;
  RECT 0.000 678.500 1.120 681.740 ;
  LAYER metal1 ;
  RECT 0.000 678.500 1.120 681.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 670.660 1.120 673.900 ;
  LAYER metal3 ;
  RECT 0.000 670.660 1.120 673.900 ;
  LAYER metal2 ;
  RECT 0.000 670.660 1.120 673.900 ;
  LAYER metal1 ;
  RECT 0.000 670.660 1.120 673.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 662.820 1.120 666.060 ;
  LAYER metal3 ;
  RECT 0.000 662.820 1.120 666.060 ;
  LAYER metal2 ;
  RECT 0.000 662.820 1.120 666.060 ;
  LAYER metal1 ;
  RECT 0.000 662.820 1.120 666.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 654.980 1.120 658.220 ;
  LAYER metal3 ;
  RECT 0.000 654.980 1.120 658.220 ;
  LAYER metal2 ;
  RECT 0.000 654.980 1.120 658.220 ;
  LAYER metal1 ;
  RECT 0.000 654.980 1.120 658.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 647.140 1.120 650.380 ;
  LAYER metal3 ;
  RECT 0.000 647.140 1.120 650.380 ;
  LAYER metal2 ;
  RECT 0.000 647.140 1.120 650.380 ;
  LAYER metal1 ;
  RECT 0.000 647.140 1.120 650.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 639.300 1.120 642.540 ;
  LAYER metal3 ;
  RECT 0.000 639.300 1.120 642.540 ;
  LAYER metal2 ;
  RECT 0.000 639.300 1.120 642.540 ;
  LAYER metal1 ;
  RECT 0.000 639.300 1.120 642.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 600.100 1.120 603.340 ;
  LAYER metal3 ;
  RECT 0.000 600.100 1.120 603.340 ;
  LAYER metal2 ;
  RECT 0.000 600.100 1.120 603.340 ;
  LAYER metal1 ;
  RECT 0.000 600.100 1.120 603.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 592.260 1.120 595.500 ;
  LAYER metal3 ;
  RECT 0.000 592.260 1.120 595.500 ;
  LAYER metal2 ;
  RECT 0.000 592.260 1.120 595.500 ;
  LAYER metal1 ;
  RECT 0.000 592.260 1.120 595.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 584.420 1.120 587.660 ;
  LAYER metal3 ;
  RECT 0.000 584.420 1.120 587.660 ;
  LAYER metal2 ;
  RECT 0.000 584.420 1.120 587.660 ;
  LAYER metal1 ;
  RECT 0.000 584.420 1.120 587.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 576.580 1.120 579.820 ;
  LAYER metal3 ;
  RECT 0.000 576.580 1.120 579.820 ;
  LAYER metal2 ;
  RECT 0.000 576.580 1.120 579.820 ;
  LAYER metal1 ;
  RECT 0.000 576.580 1.120 579.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 568.740 1.120 571.980 ;
  LAYER metal3 ;
  RECT 0.000 568.740 1.120 571.980 ;
  LAYER metal2 ;
  RECT 0.000 568.740 1.120 571.980 ;
  LAYER metal1 ;
  RECT 0.000 568.740 1.120 571.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 560.900 1.120 564.140 ;
  LAYER metal3 ;
  RECT 0.000 560.900 1.120 564.140 ;
  LAYER metal2 ;
  RECT 0.000 560.900 1.120 564.140 ;
  LAYER metal1 ;
  RECT 0.000 560.900 1.120 564.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 521.700 1.120 524.940 ;
  LAYER metal3 ;
  RECT 0.000 521.700 1.120 524.940 ;
  LAYER metal2 ;
  RECT 0.000 521.700 1.120 524.940 ;
  LAYER metal1 ;
  RECT 0.000 521.700 1.120 524.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 513.860 1.120 517.100 ;
  LAYER metal3 ;
  RECT 0.000 513.860 1.120 517.100 ;
  LAYER metal2 ;
  RECT 0.000 513.860 1.120 517.100 ;
  LAYER metal1 ;
  RECT 0.000 513.860 1.120 517.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 506.020 1.120 509.260 ;
  LAYER metal3 ;
  RECT 0.000 506.020 1.120 509.260 ;
  LAYER metal2 ;
  RECT 0.000 506.020 1.120 509.260 ;
  LAYER metal1 ;
  RECT 0.000 506.020 1.120 509.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 498.180 1.120 501.420 ;
  LAYER metal3 ;
  RECT 0.000 498.180 1.120 501.420 ;
  LAYER metal2 ;
  RECT 0.000 498.180 1.120 501.420 ;
  LAYER metal1 ;
  RECT 0.000 498.180 1.120 501.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 490.340 1.120 493.580 ;
  LAYER metal3 ;
  RECT 0.000 490.340 1.120 493.580 ;
  LAYER metal2 ;
  RECT 0.000 490.340 1.120 493.580 ;
  LAYER metal1 ;
  RECT 0.000 490.340 1.120 493.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 482.500 1.120 485.740 ;
  LAYER metal3 ;
  RECT 0.000 482.500 1.120 485.740 ;
  LAYER metal2 ;
  RECT 0.000 482.500 1.120 485.740 ;
  LAYER metal1 ;
  RECT 0.000 482.500 1.120 485.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 443.300 1.120 446.540 ;
  LAYER metal3 ;
  RECT 0.000 443.300 1.120 446.540 ;
  LAYER metal2 ;
  RECT 0.000 443.300 1.120 446.540 ;
  LAYER metal1 ;
  RECT 0.000 443.300 1.120 446.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 435.460 1.120 438.700 ;
  LAYER metal3 ;
  RECT 0.000 435.460 1.120 438.700 ;
  LAYER metal2 ;
  RECT 0.000 435.460 1.120 438.700 ;
  LAYER metal1 ;
  RECT 0.000 435.460 1.120 438.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 427.620 1.120 430.860 ;
  LAYER metal3 ;
  RECT 0.000 427.620 1.120 430.860 ;
  LAYER metal2 ;
  RECT 0.000 427.620 1.120 430.860 ;
  LAYER metal1 ;
  RECT 0.000 427.620 1.120 430.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 419.780 1.120 423.020 ;
  LAYER metal3 ;
  RECT 0.000 419.780 1.120 423.020 ;
  LAYER metal2 ;
  RECT 0.000 419.780 1.120 423.020 ;
  LAYER metal1 ;
  RECT 0.000 419.780 1.120 423.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 411.940 1.120 415.180 ;
  LAYER metal3 ;
  RECT 0.000 411.940 1.120 415.180 ;
  LAYER metal2 ;
  RECT 0.000 411.940 1.120 415.180 ;
  LAYER metal1 ;
  RECT 0.000 411.940 1.120 415.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 404.100 1.120 407.340 ;
  LAYER metal3 ;
  RECT 0.000 404.100 1.120 407.340 ;
  LAYER metal2 ;
  RECT 0.000 404.100 1.120 407.340 ;
  LAYER metal1 ;
  RECT 0.000 404.100 1.120 407.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 364.900 1.120 368.140 ;
  LAYER metal3 ;
  RECT 0.000 364.900 1.120 368.140 ;
  LAYER metal2 ;
  RECT 0.000 364.900 1.120 368.140 ;
  LAYER metal1 ;
  RECT 0.000 364.900 1.120 368.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 357.060 1.120 360.300 ;
  LAYER metal3 ;
  RECT 0.000 357.060 1.120 360.300 ;
  LAYER metal2 ;
  RECT 0.000 357.060 1.120 360.300 ;
  LAYER metal1 ;
  RECT 0.000 357.060 1.120 360.300 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 349.220 1.120 352.460 ;
  LAYER metal3 ;
  RECT 0.000 349.220 1.120 352.460 ;
  LAYER metal2 ;
  RECT 0.000 349.220 1.120 352.460 ;
  LAYER metal1 ;
  RECT 0.000 349.220 1.120 352.460 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 341.380 1.120 344.620 ;
  LAYER metal3 ;
  RECT 0.000 341.380 1.120 344.620 ;
  LAYER metal2 ;
  RECT 0.000 341.380 1.120 344.620 ;
  LAYER metal1 ;
  RECT 0.000 341.380 1.120 344.620 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 333.540 1.120 336.780 ;
  LAYER metal3 ;
  RECT 0.000 333.540 1.120 336.780 ;
  LAYER metal2 ;
  RECT 0.000 333.540 1.120 336.780 ;
  LAYER metal1 ;
  RECT 0.000 333.540 1.120 336.780 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 325.700 1.120 328.940 ;
  LAYER metal3 ;
  RECT 0.000 325.700 1.120 328.940 ;
  LAYER metal2 ;
  RECT 0.000 325.700 1.120 328.940 ;
  LAYER metal1 ;
  RECT 0.000 325.700 1.120 328.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 286.500 1.120 289.740 ;
  LAYER metal3 ;
  RECT 0.000 286.500 1.120 289.740 ;
  LAYER metal2 ;
  RECT 0.000 286.500 1.120 289.740 ;
  LAYER metal1 ;
  RECT 0.000 286.500 1.120 289.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 278.660 1.120 281.900 ;
  LAYER metal3 ;
  RECT 0.000 278.660 1.120 281.900 ;
  LAYER metal2 ;
  RECT 0.000 278.660 1.120 281.900 ;
  LAYER metal1 ;
  RECT 0.000 278.660 1.120 281.900 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 270.820 1.120 274.060 ;
  LAYER metal3 ;
  RECT 0.000 270.820 1.120 274.060 ;
  LAYER metal2 ;
  RECT 0.000 270.820 1.120 274.060 ;
  LAYER metal1 ;
  RECT 0.000 270.820 1.120 274.060 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 262.980 1.120 266.220 ;
  LAYER metal3 ;
  RECT 0.000 262.980 1.120 266.220 ;
  LAYER metal2 ;
  RECT 0.000 262.980 1.120 266.220 ;
  LAYER metal1 ;
  RECT 0.000 262.980 1.120 266.220 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 255.140 1.120 258.380 ;
  LAYER metal3 ;
  RECT 0.000 255.140 1.120 258.380 ;
  LAYER metal2 ;
  RECT 0.000 255.140 1.120 258.380 ;
  LAYER metal1 ;
  RECT 0.000 255.140 1.120 258.380 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER metal3 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER metal2 ;
  RECT 0.000 247.300 1.120 250.540 ;
  LAYER metal1 ;
  RECT 0.000 247.300 1.120 250.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER metal3 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER metal2 ;
  RECT 0.000 208.100 1.120 211.340 ;
  LAYER metal1 ;
  RECT 0.000 208.100 1.120 211.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER metal3 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER metal2 ;
  RECT 0.000 200.260 1.120 203.500 ;
  LAYER metal1 ;
  RECT 0.000 200.260 1.120 203.500 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER metal3 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER metal2 ;
  RECT 0.000 192.420 1.120 195.660 ;
  LAYER metal1 ;
  RECT 0.000 192.420 1.120 195.660 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER metal3 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER metal2 ;
  RECT 0.000 184.580 1.120 187.820 ;
  LAYER metal1 ;
  RECT 0.000 184.580 1.120 187.820 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER metal3 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER metal2 ;
  RECT 0.000 176.740 1.120 179.980 ;
  LAYER metal1 ;
  RECT 0.000 176.740 1.120 179.980 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER metal3 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER metal2 ;
  RECT 0.000 168.900 1.120 172.140 ;
  LAYER metal1 ;
  RECT 0.000 168.900 1.120 172.140 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal3 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal2 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER metal1 ;
  RECT 0.000 129.700 1.120 132.940 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal3 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal2 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER metal1 ;
  RECT 0.000 121.860 1.120 125.100 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal3 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal2 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER metal1 ;
  RECT 0.000 114.020 1.120 117.260 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal3 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal2 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER metal1 ;
  RECT 0.000 106.180 1.120 109.420 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal3 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal2 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER metal1 ;
  RECT 0.000 98.340 1.120 101.580 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal3 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal2 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER metal1 ;
  RECT 0.000 90.500 1.120 93.740 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal3 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal2 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER metal1 ;
  RECT 0.000 51.300 1.120 54.540 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal3 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal2 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER metal1 ;
  RECT 0.000 43.460 1.120 46.700 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal3 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal2 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER metal1 ;
  RECT 0.000 35.620 1.120 38.860 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal3 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal2 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER metal1 ;
  RECT 0.000 27.780 1.120 31.020 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal3 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal2 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER metal1 ;
  RECT 0.000 19.940 1.120 23.180 ;
 END
 PORT
  LAYER metal4 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal3 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal2 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER metal1 ;
  RECT 0.000 12.100 1.120 15.340 ;
 END
 PORT
  LAYER metal4 ;
  RECT 550.340 1076.880 553.880 1078.000 ;
  LAYER metal3 ;
  RECT 550.340 1076.880 553.880 1078.000 ;
  LAYER metal2 ;
  RECT 550.340 1076.880 553.880 1078.000 ;
  LAYER metal1 ;
  RECT 550.340 1076.880 553.880 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 541.660 1076.880 545.200 1078.000 ;
  LAYER metal3 ;
  RECT 541.660 1076.880 545.200 1078.000 ;
  LAYER metal2 ;
  RECT 541.660 1076.880 545.200 1078.000 ;
  LAYER metal1 ;
  RECT 541.660 1076.880 545.200 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 532.980 1076.880 536.520 1078.000 ;
  LAYER metal3 ;
  RECT 532.980 1076.880 536.520 1078.000 ;
  LAYER metal2 ;
  RECT 532.980 1076.880 536.520 1078.000 ;
  LAYER metal1 ;
  RECT 532.980 1076.880 536.520 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 489.580 1076.880 493.120 1078.000 ;
  LAYER metal3 ;
  RECT 489.580 1076.880 493.120 1078.000 ;
  LAYER metal2 ;
  RECT 489.580 1076.880 493.120 1078.000 ;
  LAYER metal1 ;
  RECT 489.580 1076.880 493.120 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 480.900 1076.880 484.440 1078.000 ;
  LAYER metal3 ;
  RECT 480.900 1076.880 484.440 1078.000 ;
  LAYER metal2 ;
  RECT 480.900 1076.880 484.440 1078.000 ;
  LAYER metal1 ;
  RECT 480.900 1076.880 484.440 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 472.220 1076.880 475.760 1078.000 ;
  LAYER metal3 ;
  RECT 472.220 1076.880 475.760 1078.000 ;
  LAYER metal2 ;
  RECT 472.220 1076.880 475.760 1078.000 ;
  LAYER metal1 ;
  RECT 472.220 1076.880 475.760 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 463.540 1076.880 467.080 1078.000 ;
  LAYER metal3 ;
  RECT 463.540 1076.880 467.080 1078.000 ;
  LAYER metal2 ;
  RECT 463.540 1076.880 467.080 1078.000 ;
  LAYER metal1 ;
  RECT 463.540 1076.880 467.080 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 454.860 1076.880 458.400 1078.000 ;
  LAYER metal3 ;
  RECT 454.860 1076.880 458.400 1078.000 ;
  LAYER metal2 ;
  RECT 454.860 1076.880 458.400 1078.000 ;
  LAYER metal1 ;
  RECT 454.860 1076.880 458.400 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 446.180 1076.880 449.720 1078.000 ;
  LAYER metal3 ;
  RECT 446.180 1076.880 449.720 1078.000 ;
  LAYER metal2 ;
  RECT 446.180 1076.880 449.720 1078.000 ;
  LAYER metal1 ;
  RECT 446.180 1076.880 449.720 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 402.780 1076.880 406.320 1078.000 ;
  LAYER metal3 ;
  RECT 402.780 1076.880 406.320 1078.000 ;
  LAYER metal2 ;
  RECT 402.780 1076.880 406.320 1078.000 ;
  LAYER metal1 ;
  RECT 402.780 1076.880 406.320 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 394.100 1076.880 397.640 1078.000 ;
  LAYER metal3 ;
  RECT 394.100 1076.880 397.640 1078.000 ;
  LAYER metal2 ;
  RECT 394.100 1076.880 397.640 1078.000 ;
  LAYER metal1 ;
  RECT 394.100 1076.880 397.640 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 385.420 1076.880 388.960 1078.000 ;
  LAYER metal3 ;
  RECT 385.420 1076.880 388.960 1078.000 ;
  LAYER metal2 ;
  RECT 385.420 1076.880 388.960 1078.000 ;
  LAYER metal1 ;
  RECT 385.420 1076.880 388.960 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 376.740 1076.880 380.280 1078.000 ;
  LAYER metal3 ;
  RECT 376.740 1076.880 380.280 1078.000 ;
  LAYER metal2 ;
  RECT 376.740 1076.880 380.280 1078.000 ;
  LAYER metal1 ;
  RECT 376.740 1076.880 380.280 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 368.060 1076.880 371.600 1078.000 ;
  LAYER metal3 ;
  RECT 368.060 1076.880 371.600 1078.000 ;
  LAYER metal2 ;
  RECT 368.060 1076.880 371.600 1078.000 ;
  LAYER metal1 ;
  RECT 368.060 1076.880 371.600 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 359.380 1076.880 362.920 1078.000 ;
  LAYER metal3 ;
  RECT 359.380 1076.880 362.920 1078.000 ;
  LAYER metal2 ;
  RECT 359.380 1076.880 362.920 1078.000 ;
  LAYER metal1 ;
  RECT 359.380 1076.880 362.920 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 315.980 1076.880 319.520 1078.000 ;
  LAYER metal3 ;
  RECT 315.980 1076.880 319.520 1078.000 ;
  LAYER metal2 ;
  RECT 315.980 1076.880 319.520 1078.000 ;
  LAYER metal1 ;
  RECT 315.980 1076.880 319.520 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 307.300 1076.880 310.840 1078.000 ;
  LAYER metal3 ;
  RECT 307.300 1076.880 310.840 1078.000 ;
  LAYER metal2 ;
  RECT 307.300 1076.880 310.840 1078.000 ;
  LAYER metal1 ;
  RECT 307.300 1076.880 310.840 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 298.620 1076.880 302.160 1078.000 ;
  LAYER metal3 ;
  RECT 298.620 1076.880 302.160 1078.000 ;
  LAYER metal2 ;
  RECT 298.620 1076.880 302.160 1078.000 ;
  LAYER metal1 ;
  RECT 298.620 1076.880 302.160 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 289.940 1076.880 293.480 1078.000 ;
  LAYER metal3 ;
  RECT 289.940 1076.880 293.480 1078.000 ;
  LAYER metal2 ;
  RECT 289.940 1076.880 293.480 1078.000 ;
  LAYER metal1 ;
  RECT 289.940 1076.880 293.480 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 281.260 1076.880 284.800 1078.000 ;
  LAYER metal3 ;
  RECT 281.260 1076.880 284.800 1078.000 ;
  LAYER metal2 ;
  RECT 281.260 1076.880 284.800 1078.000 ;
  LAYER metal1 ;
  RECT 281.260 1076.880 284.800 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 272.580 1076.880 276.120 1078.000 ;
  LAYER metal3 ;
  RECT 272.580 1076.880 276.120 1078.000 ;
  LAYER metal2 ;
  RECT 272.580 1076.880 276.120 1078.000 ;
  LAYER metal1 ;
  RECT 272.580 1076.880 276.120 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 229.180 1076.880 232.720 1078.000 ;
  LAYER metal3 ;
  RECT 229.180 1076.880 232.720 1078.000 ;
  LAYER metal2 ;
  RECT 229.180 1076.880 232.720 1078.000 ;
  LAYER metal1 ;
  RECT 229.180 1076.880 232.720 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 220.500 1076.880 224.040 1078.000 ;
  LAYER metal3 ;
  RECT 220.500 1076.880 224.040 1078.000 ;
  LAYER metal2 ;
  RECT 220.500 1076.880 224.040 1078.000 ;
  LAYER metal1 ;
  RECT 220.500 1076.880 224.040 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 211.820 1076.880 215.360 1078.000 ;
  LAYER metal3 ;
  RECT 211.820 1076.880 215.360 1078.000 ;
  LAYER metal2 ;
  RECT 211.820 1076.880 215.360 1078.000 ;
  LAYER metal1 ;
  RECT 211.820 1076.880 215.360 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 203.140 1076.880 206.680 1078.000 ;
  LAYER metal3 ;
  RECT 203.140 1076.880 206.680 1078.000 ;
  LAYER metal2 ;
  RECT 203.140 1076.880 206.680 1078.000 ;
  LAYER metal1 ;
  RECT 203.140 1076.880 206.680 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 194.460 1076.880 198.000 1078.000 ;
  LAYER metal3 ;
  RECT 194.460 1076.880 198.000 1078.000 ;
  LAYER metal2 ;
  RECT 194.460 1076.880 198.000 1078.000 ;
  LAYER metal1 ;
  RECT 194.460 1076.880 198.000 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 185.780 1076.880 189.320 1078.000 ;
  LAYER metal3 ;
  RECT 185.780 1076.880 189.320 1078.000 ;
  LAYER metal2 ;
  RECT 185.780 1076.880 189.320 1078.000 ;
  LAYER metal1 ;
  RECT 185.780 1076.880 189.320 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 142.380 1076.880 145.920 1078.000 ;
  LAYER metal3 ;
  RECT 142.380 1076.880 145.920 1078.000 ;
  LAYER metal2 ;
  RECT 142.380 1076.880 145.920 1078.000 ;
  LAYER metal1 ;
  RECT 142.380 1076.880 145.920 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 133.700 1076.880 137.240 1078.000 ;
  LAYER metal3 ;
  RECT 133.700 1076.880 137.240 1078.000 ;
  LAYER metal2 ;
  RECT 133.700 1076.880 137.240 1078.000 ;
  LAYER metal1 ;
  RECT 133.700 1076.880 137.240 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 125.020 1076.880 128.560 1078.000 ;
  LAYER metal3 ;
  RECT 125.020 1076.880 128.560 1078.000 ;
  LAYER metal2 ;
  RECT 125.020 1076.880 128.560 1078.000 ;
  LAYER metal1 ;
  RECT 125.020 1076.880 128.560 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 116.340 1076.880 119.880 1078.000 ;
  LAYER metal3 ;
  RECT 116.340 1076.880 119.880 1078.000 ;
  LAYER metal2 ;
  RECT 116.340 1076.880 119.880 1078.000 ;
  LAYER metal1 ;
  RECT 116.340 1076.880 119.880 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 107.660 1076.880 111.200 1078.000 ;
  LAYER metal3 ;
  RECT 107.660 1076.880 111.200 1078.000 ;
  LAYER metal2 ;
  RECT 107.660 1076.880 111.200 1078.000 ;
  LAYER metal1 ;
  RECT 107.660 1076.880 111.200 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 98.980 1076.880 102.520 1078.000 ;
  LAYER metal3 ;
  RECT 98.980 1076.880 102.520 1078.000 ;
  LAYER metal2 ;
  RECT 98.980 1076.880 102.520 1078.000 ;
  LAYER metal1 ;
  RECT 98.980 1076.880 102.520 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 55.580 1076.880 59.120 1078.000 ;
  LAYER metal3 ;
  RECT 55.580 1076.880 59.120 1078.000 ;
  LAYER metal2 ;
  RECT 55.580 1076.880 59.120 1078.000 ;
  LAYER metal1 ;
  RECT 55.580 1076.880 59.120 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 46.900 1076.880 50.440 1078.000 ;
  LAYER metal3 ;
  RECT 46.900 1076.880 50.440 1078.000 ;
  LAYER metal2 ;
  RECT 46.900 1076.880 50.440 1078.000 ;
  LAYER metal1 ;
  RECT 46.900 1076.880 50.440 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 38.220 1076.880 41.760 1078.000 ;
  LAYER metal3 ;
  RECT 38.220 1076.880 41.760 1078.000 ;
  LAYER metal2 ;
  RECT 38.220 1076.880 41.760 1078.000 ;
  LAYER metal1 ;
  RECT 38.220 1076.880 41.760 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 29.540 1076.880 33.080 1078.000 ;
  LAYER metal3 ;
  RECT 29.540 1076.880 33.080 1078.000 ;
  LAYER metal2 ;
  RECT 29.540 1076.880 33.080 1078.000 ;
  LAYER metal1 ;
  RECT 29.540 1076.880 33.080 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 20.860 1076.880 24.400 1078.000 ;
  LAYER metal3 ;
  RECT 20.860 1076.880 24.400 1078.000 ;
  LAYER metal2 ;
  RECT 20.860 1076.880 24.400 1078.000 ;
  LAYER metal1 ;
  RECT 20.860 1076.880 24.400 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 12.180 1076.880 15.720 1078.000 ;
  LAYER metal3 ;
  RECT 12.180 1076.880 15.720 1078.000 ;
  LAYER metal2 ;
  RECT 12.180 1076.880 15.720 1078.000 ;
  LAYER metal1 ;
  RECT 12.180 1076.880 15.720 1078.000 ;
 END
 PORT
  LAYER metal4 ;
  RECT 552.200 0.000 555.740 1.120 ;
  LAYER metal3 ;
  RECT 552.200 0.000 555.740 1.120 ;
  LAYER metal2 ;
  RECT 552.200 0.000 555.740 1.120 ;
  LAYER metal1 ;
  RECT 552.200 0.000 555.740 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 530.500 0.000 534.040 1.120 ;
  LAYER metal3 ;
  RECT 530.500 0.000 534.040 1.120 ;
  LAYER metal2 ;
  RECT 530.500 0.000 534.040 1.120 ;
  LAYER metal1 ;
  RECT 530.500 0.000 534.040 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 513.760 0.000 517.300 1.120 ;
  LAYER metal3 ;
  RECT 513.760 0.000 517.300 1.120 ;
  LAYER metal2 ;
  RECT 513.760 0.000 517.300 1.120 ;
  LAYER metal1 ;
  RECT 513.760 0.000 517.300 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 487.100 0.000 490.640 1.120 ;
  LAYER metal3 ;
  RECT 487.100 0.000 490.640 1.120 ;
  LAYER metal2 ;
  RECT 487.100 0.000 490.640 1.120 ;
  LAYER metal1 ;
  RECT 487.100 0.000 490.640 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 466.020 0.000 469.560 1.120 ;
  LAYER metal3 ;
  RECT 466.020 0.000 469.560 1.120 ;
  LAYER metal2 ;
  RECT 466.020 0.000 469.560 1.120 ;
  LAYER metal1 ;
  RECT 466.020 0.000 469.560 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 352.560 0.000 356.100 1.120 ;
  LAYER metal3 ;
  RECT 352.560 0.000 356.100 1.120 ;
  LAYER metal2 ;
  RECT 352.560 0.000 356.100 1.120 ;
  LAYER metal1 ;
  RECT 352.560 0.000 356.100 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 330.860 0.000 334.400 1.120 ;
  LAYER metal3 ;
  RECT 330.860 0.000 334.400 1.120 ;
  LAYER metal2 ;
  RECT 330.860 0.000 334.400 1.120 ;
  LAYER metal1 ;
  RECT 330.860 0.000 334.400 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 304.200 0.000 307.740 1.120 ;
  LAYER metal3 ;
  RECT 304.200 0.000 307.740 1.120 ;
  LAYER metal2 ;
  RECT 304.200 0.000 307.740 1.120 ;
  LAYER metal1 ;
  RECT 304.200 0.000 307.740 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 295.520 0.000 299.060 1.120 ;
  LAYER metal3 ;
  RECT 295.520 0.000 299.060 1.120 ;
  LAYER metal2 ;
  RECT 295.520 0.000 299.060 1.120 ;
  LAYER metal1 ;
  RECT 295.520 0.000 299.060 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 267.620 0.000 271.160 1.120 ;
  LAYER metal3 ;
  RECT 267.620 0.000 271.160 1.120 ;
  LAYER metal2 ;
  RECT 267.620 0.000 271.160 1.120 ;
  LAYER metal1 ;
  RECT 267.620 0.000 271.160 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 246.540 0.000 250.080 1.120 ;
  LAYER metal3 ;
  RECT 246.540 0.000 250.080 1.120 ;
  LAYER metal2 ;
  RECT 246.540 0.000 250.080 1.120 ;
  LAYER metal1 ;
  RECT 246.540 0.000 250.080 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER metal3 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER metal2 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER metal1 ;
  RECT 139.900 0.000 143.440 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER metal3 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER metal2 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER metal1 ;
  RECT 113.860 0.000 117.400 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER metal3 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER metal2 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER metal1 ;
  RECT 92.160 0.000 95.700 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER metal3 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER metal2 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER metal1 ;
  RECT 70.460 0.000 74.000 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER metal3 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER metal2 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER metal1 ;
  RECT 43.800 0.000 47.340 1.120 ;
 END
 PORT
  LAYER metal4 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal3 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal2 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER metal1 ;
  RECT 27.060 0.000 30.600 1.120 ;
 END
END GND
PIN DO31
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 550.000 0.000 551.120 1.120 ;
  LAYER metal3 ;
  RECT 550.000 0.000 551.120 1.120 ;
  LAYER metal2 ;
  RECT 550.000 0.000 551.120 1.120 ;
  LAYER metal1 ;
  RECT 550.000 0.000 551.120 1.120 ;
 END
END DO31
PIN DI31
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 541.320 0.000 542.440 1.120 ;
  LAYER metal3 ;
  RECT 541.320 0.000 542.440 1.120 ;
  LAYER metal2 ;
  RECT 541.320 0.000 542.440 1.120 ;
  LAYER metal1 ;
  RECT 541.320 0.000 542.440 1.120 ;
 END
END DI31
PIN DO30
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 536.980 0.000 538.100 1.120 ;
  LAYER metal3 ;
  RECT 536.980 0.000 538.100 1.120 ;
  LAYER metal2 ;
  RECT 536.980 0.000 538.100 1.120 ;
  LAYER metal1 ;
  RECT 536.980 0.000 538.100 1.120 ;
 END
END DO30
PIN DI30
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 528.300 0.000 529.420 1.120 ;
  LAYER metal3 ;
  RECT 528.300 0.000 529.420 1.120 ;
  LAYER metal2 ;
  RECT 528.300 0.000 529.420 1.120 ;
  LAYER metal1 ;
  RECT 528.300 0.000 529.420 1.120 ;
 END
END DI30
PIN DO29
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 520.240 0.000 521.360 1.120 ;
  LAYER metal3 ;
  RECT 520.240 0.000 521.360 1.120 ;
  LAYER metal2 ;
  RECT 520.240 0.000 521.360 1.120 ;
  LAYER metal1 ;
  RECT 520.240 0.000 521.360 1.120 ;
 END
END DO29
PIN DI29
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 511.560 0.000 512.680 1.120 ;
  LAYER metal3 ;
  RECT 511.560 0.000 512.680 1.120 ;
  LAYER metal2 ;
  RECT 511.560 0.000 512.680 1.120 ;
  LAYER metal1 ;
  RECT 511.560 0.000 512.680 1.120 ;
 END
END DI29
PIN DO28
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 506.600 0.000 507.720 1.120 ;
  LAYER metal3 ;
  RECT 506.600 0.000 507.720 1.120 ;
  LAYER metal2 ;
  RECT 506.600 0.000 507.720 1.120 ;
  LAYER metal1 ;
  RECT 506.600 0.000 507.720 1.120 ;
 END
END DO28
PIN DI28
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 498.540 0.000 499.660 1.120 ;
  LAYER metal3 ;
  RECT 498.540 0.000 499.660 1.120 ;
  LAYER metal2 ;
  RECT 498.540 0.000 499.660 1.120 ;
  LAYER metal1 ;
  RECT 498.540 0.000 499.660 1.120 ;
 END
END DI28
PIN DO27
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 493.580 0.000 494.700 1.120 ;
  LAYER metal3 ;
  RECT 493.580 0.000 494.700 1.120 ;
  LAYER metal2 ;
  RECT 493.580 0.000 494.700 1.120 ;
  LAYER metal1 ;
  RECT 493.580 0.000 494.700 1.120 ;
 END
END DO27
PIN DI27
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 484.900 0.000 486.020 1.120 ;
  LAYER metal3 ;
  RECT 484.900 0.000 486.020 1.120 ;
  LAYER metal2 ;
  RECT 484.900 0.000 486.020 1.120 ;
  LAYER metal1 ;
  RECT 484.900 0.000 486.020 1.120 ;
 END
END DI27
PIN DO26
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 479.940 0.000 481.060 1.120 ;
  LAYER metal3 ;
  RECT 479.940 0.000 481.060 1.120 ;
  LAYER metal2 ;
  RECT 479.940 0.000 481.060 1.120 ;
  LAYER metal1 ;
  RECT 479.940 0.000 481.060 1.120 ;
 END
END DO26
PIN DI26
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 471.880 0.000 473.000 1.120 ;
  LAYER metal3 ;
  RECT 471.880 0.000 473.000 1.120 ;
  LAYER metal2 ;
  RECT 471.880 0.000 473.000 1.120 ;
  LAYER metal1 ;
  RECT 471.880 0.000 473.000 1.120 ;
 END
END DI26
PIN DO25
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 463.820 0.000 464.940 1.120 ;
  LAYER metal3 ;
  RECT 463.820 0.000 464.940 1.120 ;
  LAYER metal2 ;
  RECT 463.820 0.000 464.940 1.120 ;
  LAYER metal1 ;
  RECT 463.820 0.000 464.940 1.120 ;
 END
END DO25
PIN DI25
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 455.140 0.000 456.260 1.120 ;
  LAYER metal3 ;
  RECT 455.140 0.000 456.260 1.120 ;
  LAYER metal2 ;
  RECT 455.140 0.000 456.260 1.120 ;
  LAYER metal1 ;
  RECT 455.140 0.000 456.260 1.120 ;
 END
END DI25
PIN DO24
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 450.180 0.000 451.300 1.120 ;
  LAYER metal3 ;
  RECT 450.180 0.000 451.300 1.120 ;
  LAYER metal2 ;
  RECT 450.180 0.000 451.300 1.120 ;
  LAYER metal1 ;
  RECT 450.180 0.000 451.300 1.120 ;
 END
END DO24
PIN DI24
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 442.120 0.000 443.240 1.120 ;
  LAYER metal3 ;
  RECT 442.120 0.000 443.240 1.120 ;
  LAYER metal2 ;
  RECT 442.120 0.000 443.240 1.120 ;
  LAYER metal1 ;
  RECT 442.120 0.000 443.240 1.120 ;
 END
END DI24
PIN DO23
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 437.160 0.000 438.280 1.120 ;
  LAYER metal3 ;
  RECT 437.160 0.000 438.280 1.120 ;
  LAYER metal2 ;
  RECT 437.160 0.000 438.280 1.120 ;
  LAYER metal1 ;
  RECT 437.160 0.000 438.280 1.120 ;
 END
END DO23
PIN DI23
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 428.480 0.000 429.600 1.120 ;
  LAYER metal3 ;
  RECT 428.480 0.000 429.600 1.120 ;
  LAYER metal2 ;
  RECT 428.480 0.000 429.600 1.120 ;
  LAYER metal1 ;
  RECT 428.480 0.000 429.600 1.120 ;
 END
END DI23
PIN DO22
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 423.520 0.000 424.640 1.120 ;
  LAYER metal3 ;
  RECT 423.520 0.000 424.640 1.120 ;
  LAYER metal2 ;
  RECT 423.520 0.000 424.640 1.120 ;
  LAYER metal1 ;
  RECT 423.520 0.000 424.640 1.120 ;
 END
END DO22
PIN DI22
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 415.460 0.000 416.580 1.120 ;
  LAYER metal3 ;
  RECT 415.460 0.000 416.580 1.120 ;
  LAYER metal2 ;
  RECT 415.460 0.000 416.580 1.120 ;
  LAYER metal1 ;
  RECT 415.460 0.000 416.580 1.120 ;
 END
END DI22
PIN DO21
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 406.780 0.000 407.900 1.120 ;
  LAYER metal3 ;
  RECT 406.780 0.000 407.900 1.120 ;
  LAYER metal2 ;
  RECT 406.780 0.000 407.900 1.120 ;
  LAYER metal1 ;
  RECT 406.780 0.000 407.900 1.120 ;
 END
END DO21
PIN DI21
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 398.720 0.000 399.840 1.120 ;
  LAYER metal3 ;
  RECT 398.720 0.000 399.840 1.120 ;
  LAYER metal2 ;
  RECT 398.720 0.000 399.840 1.120 ;
  LAYER metal1 ;
  RECT 398.720 0.000 399.840 1.120 ;
 END
END DI21
PIN DO20
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 393.760 0.000 394.880 1.120 ;
  LAYER metal3 ;
  RECT 393.760 0.000 394.880 1.120 ;
  LAYER metal2 ;
  RECT 393.760 0.000 394.880 1.120 ;
  LAYER metal1 ;
  RECT 393.760 0.000 394.880 1.120 ;
 END
END DO20
PIN DI20
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 385.080 0.000 386.200 1.120 ;
  LAYER metal3 ;
  RECT 385.080 0.000 386.200 1.120 ;
  LAYER metal2 ;
  RECT 385.080 0.000 386.200 1.120 ;
  LAYER metal1 ;
  RECT 385.080 0.000 386.200 1.120 ;
 END
END DI20
PIN DO19
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 380.740 0.000 381.860 1.120 ;
  LAYER metal3 ;
  RECT 380.740 0.000 381.860 1.120 ;
  LAYER metal2 ;
  RECT 380.740 0.000 381.860 1.120 ;
  LAYER metal1 ;
  RECT 380.740 0.000 381.860 1.120 ;
 END
END DO19
PIN DI19
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 372.060 0.000 373.180 1.120 ;
  LAYER metal3 ;
  RECT 372.060 0.000 373.180 1.120 ;
  LAYER metal2 ;
  RECT 372.060 0.000 373.180 1.120 ;
  LAYER metal1 ;
  RECT 372.060 0.000 373.180 1.120 ;
 END
END DI19
PIN DO18
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 367.100 0.000 368.220 1.120 ;
  LAYER metal3 ;
  RECT 367.100 0.000 368.220 1.120 ;
  LAYER metal2 ;
  RECT 367.100 0.000 368.220 1.120 ;
  LAYER metal1 ;
  RECT 367.100 0.000 368.220 1.120 ;
 END
END DO18
PIN DI18
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER metal3 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER metal2 ;
  RECT 359.040 0.000 360.160 1.120 ;
  LAYER metal1 ;
  RECT 359.040 0.000 360.160 1.120 ;
 END
END DI18
PIN DO17
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 350.360 0.000 351.480 1.120 ;
  LAYER metal3 ;
  RECT 350.360 0.000 351.480 1.120 ;
  LAYER metal2 ;
  RECT 350.360 0.000 351.480 1.120 ;
  LAYER metal1 ;
  RECT 350.360 0.000 351.480 1.120 ;
 END
END DO17
PIN DI17
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 342.300 0.000 343.420 1.120 ;
  LAYER metal3 ;
  RECT 342.300 0.000 343.420 1.120 ;
  LAYER metal2 ;
  RECT 342.300 0.000 343.420 1.120 ;
  LAYER metal1 ;
  RECT 342.300 0.000 343.420 1.120 ;
 END
END DI17
PIN DO16
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 337.340 0.000 338.460 1.120 ;
  LAYER metal3 ;
  RECT 337.340 0.000 338.460 1.120 ;
  LAYER metal2 ;
  RECT 337.340 0.000 338.460 1.120 ;
  LAYER metal1 ;
  RECT 337.340 0.000 338.460 1.120 ;
 END
END DO16
PIN DI16
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 328.660 0.000 329.780 1.120 ;
  LAYER metal3 ;
  RECT 328.660 0.000 329.780 1.120 ;
  LAYER metal2 ;
  RECT 328.660 0.000 329.780 1.120 ;
  LAYER metal1 ;
  RECT 328.660 0.000 329.780 1.120 ;
 END
END DI16
PIN A1
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 323.080 0.000 324.200 1.120 ;
  LAYER metal3 ;
  RECT 323.080 0.000 324.200 1.120 ;
  LAYER metal2 ;
  RECT 323.080 0.000 324.200 1.120 ;
  LAYER metal1 ;
  RECT 323.080 0.000 324.200 1.120 ;
 END
END A1
PIN WEB
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER metal4 ;
  RECT 321.220 0.000 322.340 1.120 ;
  LAYER metal3 ;
  RECT 321.220 0.000 322.340 1.120 ;
  LAYER metal2 ;
  RECT 321.220 0.000 322.340 1.120 ;
  LAYER metal1 ;
  RECT 321.220 0.000 322.340 1.120 ;
 END
END WEB
PIN OE
  DIRECTION INPUT ;
  CAPACITANCE 0.033 ;
 PORT
  LAYER metal4 ;
  RECT 316.260 0.000 317.380 1.120 ;
  LAYER metal3 ;
  RECT 316.260 0.000 317.380 1.120 ;
  LAYER metal2 ;
  RECT 316.260 0.000 317.380 1.120 ;
  LAYER metal1 ;
  RECT 316.260 0.000 317.380 1.120 ;
 END
END OE
PIN CS
  DIRECTION INPUT ;
  CAPACITANCE 0.123 ;
 PORT
  LAYER metal4 ;
  RECT 314.400 0.000 315.520 1.120 ;
  LAYER metal3 ;
  RECT 314.400 0.000 315.520 1.120 ;
  LAYER metal2 ;
  RECT 314.400 0.000 315.520 1.120 ;
  LAYER metal1 ;
  RECT 314.400 0.000 315.520 1.120 ;
 END
END CS
PIN A2
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 293.320 0.000 294.440 1.120 ;
  LAYER metal3 ;
  RECT 293.320 0.000 294.440 1.120 ;
  LAYER metal2 ;
  RECT 293.320 0.000 294.440 1.120 ;
  LAYER metal1 ;
  RECT 293.320 0.000 294.440 1.120 ;
 END
END A2
PIN CK
  DIRECTION INPUT ;
  CAPACITANCE 0.063 ;
 PORT
  LAYER metal4 ;
  RECT 290.220 0.000 291.340 1.120 ;
  LAYER metal3 ;
  RECT 290.220 0.000 291.340 1.120 ;
  LAYER metal2 ;
  RECT 290.220 0.000 291.340 1.120 ;
  LAYER metal1 ;
  RECT 290.220 0.000 291.340 1.120 ;
 END
END CK
PIN A0
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 287.740 0.000 288.860 1.120 ;
  LAYER metal3 ;
  RECT 287.740 0.000 288.860 1.120 ;
  LAYER metal2 ;
  RECT 287.740 0.000 288.860 1.120 ;
  LAYER metal1 ;
  RECT 287.740 0.000 288.860 1.120 ;
 END
END A0
PIN A3
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 283.400 0.000 284.520 1.120 ;
  LAYER metal3 ;
  RECT 283.400 0.000 284.520 1.120 ;
  LAYER metal2 ;
  RECT 283.400 0.000 284.520 1.120 ;
  LAYER metal1 ;
  RECT 283.400 0.000 284.520 1.120 ;
 END
END A3
PIN A4
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 275.960 0.000 277.080 1.120 ;
  LAYER metal3 ;
  RECT 275.960 0.000 277.080 1.120 ;
  LAYER metal2 ;
  RECT 275.960 0.000 277.080 1.120 ;
  LAYER metal1 ;
  RECT 275.960 0.000 277.080 1.120 ;
 END
END A4
PIN A5
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 272.860 0.000 273.980 1.120 ;
  LAYER metal3 ;
  RECT 272.860 0.000 273.980 1.120 ;
  LAYER metal2 ;
  RECT 272.860 0.000 273.980 1.120 ;
  LAYER metal1 ;
  RECT 272.860 0.000 273.980 1.120 ;
 END
END A5
PIN A6
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 265.420 0.000 266.540 1.120 ;
  LAYER metal3 ;
  RECT 265.420 0.000 266.540 1.120 ;
  LAYER metal2 ;
  RECT 265.420 0.000 266.540 1.120 ;
  LAYER metal1 ;
  RECT 265.420 0.000 266.540 1.120 ;
 END
END A6
PIN A7
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 262.320 0.000 263.440 1.120 ;
  LAYER metal3 ;
  RECT 262.320 0.000 263.440 1.120 ;
  LAYER metal2 ;
  RECT 262.320 0.000 263.440 1.120 ;
  LAYER metal1 ;
  RECT 262.320 0.000 263.440 1.120 ;
 END
END A7
PIN A8
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER metal3 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER metal2 ;
  RECT 254.880 0.000 256.000 1.120 ;
  LAYER metal1 ;
  RECT 254.880 0.000 256.000 1.120 ;
 END
END A8
PIN A9
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 251.780 0.000 252.900 1.120 ;
  LAYER metal3 ;
  RECT 251.780 0.000 252.900 1.120 ;
  LAYER metal2 ;
  RECT 251.780 0.000 252.900 1.120 ;
  LAYER metal1 ;
  RECT 251.780 0.000 252.900 1.120 ;
 END
END A9
PIN A10
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 244.340 0.000 245.460 1.120 ;
  LAYER metal3 ;
  RECT 244.340 0.000 245.460 1.120 ;
  LAYER metal2 ;
  RECT 244.340 0.000 245.460 1.120 ;
  LAYER metal1 ;
  RECT 244.340 0.000 245.460 1.120 ;
 END
END A10
PIN A11
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER metal4 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER metal3 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER metal2 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER metal1 ;
  RECT 241.240 0.000 242.360 1.120 ;
 END
END A11
PIN DO15
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER metal3 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER metal2 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER metal1 ;
  RECT 233.180 0.000 234.300 1.120 ;
 END
END DO15
PIN DI15
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER metal3 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER metal2 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER metal1 ;
  RECT 224.500 0.000 225.620 1.120 ;
 END
END DI15
PIN DO14
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER metal3 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER metal2 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER metal1 ;
  RECT 219.540 0.000 220.660 1.120 ;
 END
END DO14
PIN DI14
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER metal3 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER metal2 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER metal1 ;
  RECT 211.480 0.000 212.600 1.120 ;
 END
END DI14
PIN DO13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER metal3 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER metal2 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER metal1 ;
  RECT 202.800 0.000 203.920 1.120 ;
 END
END DO13
PIN DI13
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER metal3 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER metal2 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER metal1 ;
  RECT 194.740 0.000 195.860 1.120 ;
 END
END DI13
PIN DO12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER metal3 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER metal2 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER metal1 ;
  RECT 189.780 0.000 190.900 1.120 ;
 END
END DO12
PIN DI12
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER metal3 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER metal2 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER metal1 ;
  RECT 181.100 0.000 182.220 1.120 ;
 END
END DI12
PIN DO11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER metal3 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER metal2 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER metal1 ;
  RECT 176.140 0.000 177.260 1.120 ;
 END
END DO11
PIN DI11
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER metal3 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER metal2 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER metal1 ;
  RECT 168.080 0.000 169.200 1.120 ;
 END
END DI11
PIN DO10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER metal3 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER metal2 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER metal1 ;
  RECT 163.120 0.000 164.240 1.120 ;
 END
END DO10
PIN DI10
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER metal3 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER metal2 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER metal1 ;
  RECT 154.440 0.000 155.560 1.120 ;
 END
END DI10
PIN DO9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER metal3 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER metal2 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER metal1 ;
  RECT 146.380 0.000 147.500 1.120 ;
 END
END DO9
PIN DI9
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER metal3 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER metal2 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER metal1 ;
  RECT 137.700 0.000 138.820 1.120 ;
 END
END DI9
PIN DO8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER metal3 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER metal2 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER metal1 ;
  RECT 133.360 0.000 134.480 1.120 ;
 END
END DO8
PIN DI8
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER metal3 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER metal2 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER metal1 ;
  RECT 124.680 0.000 125.800 1.120 ;
 END
END DI8
PIN DO7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER metal3 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER metal2 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER metal1 ;
  RECT 119.720 0.000 120.840 1.120 ;
 END
END DO7
PIN DI7
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER metal3 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER metal2 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER metal1 ;
  RECT 111.660 0.000 112.780 1.120 ;
 END
END DI7
PIN DO6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal3 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal2 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER metal1 ;
  RECT 106.700 0.000 107.820 1.120 ;
 END
END DO6
PIN DI6
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER metal3 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER metal2 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER metal1 ;
  RECT 98.020 0.000 99.140 1.120 ;
 END
END DI6
PIN DO5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER metal3 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER metal2 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER metal1 ;
  RECT 89.960 0.000 91.080 1.120 ;
 END
END DO5
PIN DI5
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER metal3 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER metal2 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER metal1 ;
  RECT 81.280 0.000 82.400 1.120 ;
 END
END DI5
PIN DO4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER metal3 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER metal2 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER metal1 ;
  RECT 76.320 0.000 77.440 1.120 ;
 END
END DO4
PIN DI4
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER metal3 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER metal2 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER metal1 ;
  RECT 68.260 0.000 69.380 1.120 ;
 END
END DI4
PIN DO3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER metal3 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER metal2 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER metal1 ;
  RECT 63.300 0.000 64.420 1.120 ;
 END
END DO3
PIN DI3
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER metal3 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER metal2 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER metal1 ;
  RECT 54.620 0.000 55.740 1.120 ;
 END
END DI3
PIN DO2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER metal3 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER metal2 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER metal1 ;
  RECT 50.280 0.000 51.400 1.120 ;
 END
END DO2
PIN DI2
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER metal3 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER metal2 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER metal1 ;
  RECT 41.600 0.000 42.720 1.120 ;
 END
END DI2
PIN DO1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal3 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal2 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER metal1 ;
  RECT 33.540 0.000 34.660 1.120 ;
 END
END DO1
PIN DI1
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal3 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal2 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER metal1 ;
  RECT 24.860 0.000 25.980 1.120 ;
 END
END DI1
PIN DO0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER metal4 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal3 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal2 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER metal1 ;
  RECT 19.900 0.000 21.020 1.120 ;
 END
END DO0
PIN DI0
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER metal4 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal3 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal2 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER metal1 ;
  RECT 11.840 0.000 12.960 1.120 ;
 END
END DI0
OBS
  LAYER metal1 SPACING 0.280 ;
  RECT 0.000 0.140 563.580 1078.000 ;
  LAYER metal2 SPACING 0.320 ;
  RECT 0.000 0.140 563.580 1078.000 ;
  LAYER metal3 SPACING 0.320 ;
  RECT 0.000 0.140 563.580 1078.000 ;
  LAYER metal4 SPACING 0.600 ;
  RECT 0.000 0.140 563.580 1078.000 ;
  LAYER via ;
  RECT 0.000 0.140 563.580 1078.000 ;
  LAYER via2 ;
  RECT 0.000 0.140 563.580 1078.000 ;
  LAYER via3 ;
  RECT 0.000 0.140 563.580 1078.000 ;
END
END dma_sram
END LIBRARY



